package data_types; endpackage