
module adder_full(a,b,cin,cout,s);
input a,b,cin;
output s,cout;
wire r,r1,r2;
xor(s,a,b,cin);
and(r,a,b);
and(r1,b,cin);
and(r2,a,cin);
or(cout,r,r1,r2);
endmodule

module adder_half(input a,input b,output cout,output s);
xor(s,a,b);
and(cout,a,b);
endmodule

module dadda(input [31:0]a,input [31:0]b,output [63:0]p);

wire [31:0]pr_and1;

wire [31:0]pr_and2;

wire [31:0]pr_and3;

wire [31:0]pr_and4;

wire [31:0]pr_and5;

wire [31:0]pr_and6;

wire [31:0]pr_and7;

wire [31:0]pr_and8;

wire [31:0]pr_and9;

wire [31:0]pr_and10;

wire [31:0]pr_and11;

wire [31:0]pr_and12;

wire [31:0]pr_and13;

wire [31:0]pr_and14;

wire [31:0]pr_and15;

wire [31:0]pr_and16;

wire [31:0]pr_and17;

wire [31:0]pr_and18;

wire [31:0]pr_and19;

wire [31:0]pr_and20;

wire [31:0]pr_and21;

wire [31:0]pr_and22;

wire [31:0]pr_and23;

wire [31:0]pr_and24;

wire [31:0]pr_and25;

wire [31:0]pr_and26;

wire [31:0]pr_and27;

wire [31:0]pr_and28;

wire [31:0]pr_and29;

wire [31:0]pr_and30;

wire [31:0]pr_and31;

wire [31:0]pr_and32;


wire [30:0]s1;
wire [31:0]c1;

wire [30:0]s2;
wire [31:0]c2;

wire [30:0]s3;
wire [31:0]c3;

wire [30:0]s4;
wire [31:0]c4;

wire [30:0]s5;
wire [31:0]c5;

wire [30:0]s6;
wire [31:0]c6;

wire [30:0]s7;
wire [31:0]c7;

wire [30:0]s8;
wire [31:0]c8;

wire [30:0]s9;
wire [31:0]c9;

wire [30:0]s10;
wire [31:0]c10;

wire [30:0]s11;
wire [31:0]c11;

wire [30:0]s12;
wire [31:0]c12;

wire [30:0]s13;
wire [31:0]c13;

wire [30:0]s14;
wire [31:0]c14;

wire [30:0]s15;
wire [31:0]c15;

wire [30:0]s16;
wire [31:0]c16;

wire [30:0]s17;
wire [31:0]c17;

wire [30:0]s18;
wire [31:0]c18;

wire [30:0]s19;
wire [31:0]c19;

wire [30:0]s20;
wire [31:0]c20;

wire [30:0]s21;
wire [31:0]c21;

wire [30:0]s22;
wire [31:0]c22;

wire [30:0]s23;
wire [31:0]c23;

wire [30:0]s24;
wire [31:0]c24;

wire [30:0]s25;
wire [31:0]c25;

wire [30:0]s26;
wire [31:0]c26;

wire [30:0]s27;
wire [31:0]c27;

wire [30:0]s28;
wire [31:0]c28;

wire [30:0]s29;
wire [31:0]c29;

wire [30:0]s30;
wire [31:0]c30;

wire [31:0]c31;
wire c;
// wire [63:0]p;
wire [31:0]si;



        and(pr_and1[0],b[0],a[0]);


        and(pr_and1[1],b[0],a[1]);


        and(pr_and1[2],b[0],a[2]);


        and(pr_and1[3],b[0],a[3]);


        and(pr_and1[4],b[0],a[4]);


        and(pr_and1[5],b[0],a[5]);


        and(pr_and1[6],b[0],a[6]);


        and(pr_and1[7],b[0],a[7]);


        and(pr_and1[8],b[0],a[8]);


        and(pr_and1[9],b[0],a[9]);


        and(pr_and1[10],b[0],a[10]);


        and(pr_and1[11],b[0],a[11]);


        and(pr_and1[12],b[0],a[12]);


        and(pr_and1[13],b[0],a[13]);


        and(pr_and1[14],b[0],a[14]);


        and(pr_and1[15],b[0],a[15]);


        and(pr_and1[16],b[0],a[16]);


        and(pr_and1[17],b[0],a[17]);


        and(pr_and1[18],b[0],a[18]);


        and(pr_and1[19],b[0],a[19]);


        and(pr_and1[20],b[0],a[20]);


        and(pr_and1[21],b[0],a[21]);


        and(pr_and1[22],b[0],a[22]);


        and(pr_and1[23],b[0],a[23]);


        and(pr_and1[24],b[0],a[24]);


        and(pr_and1[25],b[0],a[25]);


        and(pr_and1[26],b[0],a[26]);


        and(pr_and1[27],b[0],a[27]);


        and(pr_and1[28],b[0],a[28]);


        and(pr_and1[29],b[0],a[29]);


        and(pr_and1[30],b[0],a[30]);


        and(pr_and1[31],b[0],a[31]);


    not(si[0],pr_and1[31]);


        and(pr_and2[0],b[1],a[0]);


        and(pr_and2[1],b[1],a[1]);


        and(pr_and2[2],b[1],a[2]);


        and(pr_and2[3],b[1],a[3]);


        and(pr_and2[4],b[1],a[4]);


        and(pr_and2[5],b[1],a[5]);


        and(pr_and2[6],b[1],a[6]);


        and(pr_and2[7],b[1],a[7]);


        and(pr_and2[8],b[1],a[8]);


        and(pr_and2[9],b[1],a[9]);


        and(pr_and2[10],b[1],a[10]);


        and(pr_and2[11],b[1],a[11]);


        and(pr_and2[12],b[1],a[12]);


        and(pr_and2[13],b[1],a[13]);


        and(pr_and2[14],b[1],a[14]);


        and(pr_and2[15],b[1],a[15]);


        and(pr_and2[16],b[1],a[16]);


        and(pr_and2[17],b[1],a[17]);


        and(pr_and2[18],b[1],a[18]);


        and(pr_and2[19],b[1],a[19]);


        and(pr_and2[20],b[1],a[20]);


        and(pr_and2[21],b[1],a[21]);


        and(pr_and2[22],b[1],a[22]);


        and(pr_and2[23],b[1],a[23]);


        and(pr_and2[24],b[1],a[24]);


        and(pr_and2[25],b[1],a[25]);


        and(pr_and2[26],b[1],a[26]);


        and(pr_and2[27],b[1],a[27]);


        and(pr_and2[28],b[1],a[28]);


        and(pr_and2[29],b[1],a[29]);


        and(pr_and2[30],b[1],a[30]);


        and(pr_and2[31],b[1],a[31]);


    not(si[1],pr_and2[31]);


        and(pr_and3[0],b[2],a[0]);


        and(pr_and3[1],b[2],a[1]);


        and(pr_and3[2],b[2],a[2]);


        and(pr_and3[3],b[2],a[3]);


        and(pr_and3[4],b[2],a[4]);


        and(pr_and3[5],b[2],a[5]);


        and(pr_and3[6],b[2],a[6]);


        and(pr_and3[7],b[2],a[7]);


        and(pr_and3[8],b[2],a[8]);


        and(pr_and3[9],b[2],a[9]);


        and(pr_and3[10],b[2],a[10]);


        and(pr_and3[11],b[2],a[11]);


        and(pr_and3[12],b[2],a[12]);


        and(pr_and3[13],b[2],a[13]);


        and(pr_and3[14],b[2],a[14]);


        and(pr_and3[15],b[2],a[15]);


        and(pr_and3[16],b[2],a[16]);


        and(pr_and3[17],b[2],a[17]);


        and(pr_and3[18],b[2],a[18]);


        and(pr_and3[19],b[2],a[19]);


        and(pr_and3[20],b[2],a[20]);


        and(pr_and3[21],b[2],a[21]);


        and(pr_and3[22],b[2],a[22]);


        and(pr_and3[23],b[2],a[23]);


        and(pr_and3[24],b[2],a[24]);


        and(pr_and3[25],b[2],a[25]);


        and(pr_and3[26],b[2],a[26]);


        and(pr_and3[27],b[2],a[27]);


        and(pr_and3[28],b[2],a[28]);


        and(pr_and3[29],b[2],a[29]);


        and(pr_and3[30],b[2],a[30]);


        and(pr_and3[31],b[2],a[31]);


    not(si[2],pr_and3[31]);


        and(pr_and4[0],b[3],a[0]);


        and(pr_and4[1],b[3],a[1]);


        and(pr_and4[2],b[3],a[2]);


        and(pr_and4[3],b[3],a[3]);


        and(pr_and4[4],b[3],a[4]);


        and(pr_and4[5],b[3],a[5]);


        and(pr_and4[6],b[3],a[6]);


        and(pr_and4[7],b[3],a[7]);


        and(pr_and4[8],b[3],a[8]);


        and(pr_and4[9],b[3],a[9]);


        and(pr_and4[10],b[3],a[10]);


        and(pr_and4[11],b[3],a[11]);


        and(pr_and4[12],b[3],a[12]);


        and(pr_and4[13],b[3],a[13]);


        and(pr_and4[14],b[3],a[14]);


        and(pr_and4[15],b[3],a[15]);


        and(pr_and4[16],b[3],a[16]);


        and(pr_and4[17],b[3],a[17]);


        and(pr_and4[18],b[3],a[18]);


        and(pr_and4[19],b[3],a[19]);


        and(pr_and4[20],b[3],a[20]);


        and(pr_and4[21],b[3],a[21]);


        and(pr_and4[22],b[3],a[22]);


        and(pr_and4[23],b[3],a[23]);


        and(pr_and4[24],b[3],a[24]);


        and(pr_and4[25],b[3],a[25]);


        and(pr_and4[26],b[3],a[26]);


        and(pr_and4[27],b[3],a[27]);


        and(pr_and4[28],b[3],a[28]);


        and(pr_and4[29],b[3],a[29]);


        and(pr_and4[30],b[3],a[30]);


        and(pr_and4[31],b[3],a[31]);


    not(si[3],pr_and4[31]);


        and(pr_and5[0],b[4],a[0]);


        and(pr_and5[1],b[4],a[1]);


        and(pr_and5[2],b[4],a[2]);


        and(pr_and5[3],b[4],a[3]);


        and(pr_and5[4],b[4],a[4]);


        and(pr_and5[5],b[4],a[5]);


        and(pr_and5[6],b[4],a[6]);


        and(pr_and5[7],b[4],a[7]);


        and(pr_and5[8],b[4],a[8]);


        and(pr_and5[9],b[4],a[9]);


        and(pr_and5[10],b[4],a[10]);


        and(pr_and5[11],b[4],a[11]);


        and(pr_and5[12],b[4],a[12]);


        and(pr_and5[13],b[4],a[13]);


        and(pr_and5[14],b[4],a[14]);


        and(pr_and5[15],b[4],a[15]);


        and(pr_and5[16],b[4],a[16]);


        and(pr_and5[17],b[4],a[17]);


        and(pr_and5[18],b[4],a[18]);


        and(pr_and5[19],b[4],a[19]);


        and(pr_and5[20],b[4],a[20]);


        and(pr_and5[21],b[4],a[21]);


        and(pr_and5[22],b[4],a[22]);


        and(pr_and5[23],b[4],a[23]);


        and(pr_and5[24],b[4],a[24]);


        and(pr_and5[25],b[4],a[25]);


        and(pr_and5[26],b[4],a[26]);


        and(pr_and5[27],b[4],a[27]);


        and(pr_and5[28],b[4],a[28]);


        and(pr_and5[29],b[4],a[29]);


        and(pr_and5[30],b[4],a[30]);


        and(pr_and5[31],b[4],a[31]);


    not(si[4],pr_and5[31]);


        and(pr_and6[0],b[5],a[0]);


        and(pr_and6[1],b[5],a[1]);


        and(pr_and6[2],b[5],a[2]);


        and(pr_and6[3],b[5],a[3]);


        and(pr_and6[4],b[5],a[4]);


        and(pr_and6[5],b[5],a[5]);


        and(pr_and6[6],b[5],a[6]);


        and(pr_and6[7],b[5],a[7]);


        and(pr_and6[8],b[5],a[8]);


        and(pr_and6[9],b[5],a[9]);


        and(pr_and6[10],b[5],a[10]);


        and(pr_and6[11],b[5],a[11]);


        and(pr_and6[12],b[5],a[12]);


        and(pr_and6[13],b[5],a[13]);


        and(pr_and6[14],b[5],a[14]);


        and(pr_and6[15],b[5],a[15]);


        and(pr_and6[16],b[5],a[16]);


        and(pr_and6[17],b[5],a[17]);


        and(pr_and6[18],b[5],a[18]);


        and(pr_and6[19],b[5],a[19]);


        and(pr_and6[20],b[5],a[20]);


        and(pr_and6[21],b[5],a[21]);


        and(pr_and6[22],b[5],a[22]);


        and(pr_and6[23],b[5],a[23]);


        and(pr_and6[24],b[5],a[24]);


        and(pr_and6[25],b[5],a[25]);


        and(pr_and6[26],b[5],a[26]);


        and(pr_and6[27],b[5],a[27]);


        and(pr_and6[28],b[5],a[28]);


        and(pr_and6[29],b[5],a[29]);


        and(pr_and6[30],b[5],a[30]);


        and(pr_and6[31],b[5],a[31]);


    not(si[5],pr_and6[31]);


        and(pr_and7[0],b[6],a[0]);


        and(pr_and7[1],b[6],a[1]);


        and(pr_and7[2],b[6],a[2]);


        and(pr_and7[3],b[6],a[3]);


        and(pr_and7[4],b[6],a[4]);


        and(pr_and7[5],b[6],a[5]);


        and(pr_and7[6],b[6],a[6]);


        and(pr_and7[7],b[6],a[7]);


        and(pr_and7[8],b[6],a[8]);


        and(pr_and7[9],b[6],a[9]);


        and(pr_and7[10],b[6],a[10]);


        and(pr_and7[11],b[6],a[11]);


        and(pr_and7[12],b[6],a[12]);


        and(pr_and7[13],b[6],a[13]);


        and(pr_and7[14],b[6],a[14]);


        and(pr_and7[15],b[6],a[15]);


        and(pr_and7[16],b[6],a[16]);


        and(pr_and7[17],b[6],a[17]);


        and(pr_and7[18],b[6],a[18]);


        and(pr_and7[19],b[6],a[19]);


        and(pr_and7[20],b[6],a[20]);


        and(pr_and7[21],b[6],a[21]);


        and(pr_and7[22],b[6],a[22]);


        and(pr_and7[23],b[6],a[23]);


        and(pr_and7[24],b[6],a[24]);


        and(pr_and7[25],b[6],a[25]);


        and(pr_and7[26],b[6],a[26]);


        and(pr_and7[27],b[6],a[27]);


        and(pr_and7[28],b[6],a[28]);


        and(pr_and7[29],b[6],a[29]);


        and(pr_and7[30],b[6],a[30]);


        and(pr_and7[31],b[6],a[31]);


    not(si[6],pr_and7[31]);


        and(pr_and8[0],b[7],a[0]);


        and(pr_and8[1],b[7],a[1]);


        and(pr_and8[2],b[7],a[2]);


        and(pr_and8[3],b[7],a[3]);


        and(pr_and8[4],b[7],a[4]);


        and(pr_and8[5],b[7],a[5]);


        and(pr_and8[6],b[7],a[6]);


        and(pr_and8[7],b[7],a[7]);


        and(pr_and8[8],b[7],a[8]);


        and(pr_and8[9],b[7],a[9]);


        and(pr_and8[10],b[7],a[10]);


        and(pr_and8[11],b[7],a[11]);


        and(pr_and8[12],b[7],a[12]);


        and(pr_and8[13],b[7],a[13]);


        and(pr_and8[14],b[7],a[14]);


        and(pr_and8[15],b[7],a[15]);


        and(pr_and8[16],b[7],a[16]);


        and(pr_and8[17],b[7],a[17]);


        and(pr_and8[18],b[7],a[18]);


        and(pr_and8[19],b[7],a[19]);


        and(pr_and8[20],b[7],a[20]);


        and(pr_and8[21],b[7],a[21]);


        and(pr_and8[22],b[7],a[22]);


        and(pr_and8[23],b[7],a[23]);


        and(pr_and8[24],b[7],a[24]);


        and(pr_and8[25],b[7],a[25]);


        and(pr_and8[26],b[7],a[26]);


        and(pr_and8[27],b[7],a[27]);


        and(pr_and8[28],b[7],a[28]);


        and(pr_and8[29],b[7],a[29]);


        and(pr_and8[30],b[7],a[30]);


        and(pr_and8[31],b[7],a[31]);


    not(si[7],pr_and8[31]);


        and(pr_and9[0],b[8],a[0]);


        and(pr_and9[1],b[8],a[1]);


        and(pr_and9[2],b[8],a[2]);


        and(pr_and9[3],b[8],a[3]);


        and(pr_and9[4],b[8],a[4]);


        and(pr_and9[5],b[8],a[5]);


        and(pr_and9[6],b[8],a[6]);


        and(pr_and9[7],b[8],a[7]);


        and(pr_and9[8],b[8],a[8]);


        and(pr_and9[9],b[8],a[9]);


        and(pr_and9[10],b[8],a[10]);


        and(pr_and9[11],b[8],a[11]);


        and(pr_and9[12],b[8],a[12]);


        and(pr_and9[13],b[8],a[13]);


        and(pr_and9[14],b[8],a[14]);


        and(pr_and9[15],b[8],a[15]);


        and(pr_and9[16],b[8],a[16]);


        and(pr_and9[17],b[8],a[17]);


        and(pr_and9[18],b[8],a[18]);


        and(pr_and9[19],b[8],a[19]);


        and(pr_and9[20],b[8],a[20]);


        and(pr_and9[21],b[8],a[21]);


        and(pr_and9[22],b[8],a[22]);


        and(pr_and9[23],b[8],a[23]);


        and(pr_and9[24],b[8],a[24]);


        and(pr_and9[25],b[8],a[25]);


        and(pr_and9[26],b[8],a[26]);


        and(pr_and9[27],b[8],a[27]);


        and(pr_and9[28],b[8],a[28]);


        and(pr_and9[29],b[8],a[29]);


        and(pr_and9[30],b[8],a[30]);


        and(pr_and9[31],b[8],a[31]);


    not(si[8],pr_and9[31]);


        and(pr_and10[0],b[9],a[0]);


        and(pr_and10[1],b[9],a[1]);


        and(pr_and10[2],b[9],a[2]);


        and(pr_and10[3],b[9],a[3]);


        and(pr_and10[4],b[9],a[4]);


        and(pr_and10[5],b[9],a[5]);


        and(pr_and10[6],b[9],a[6]);


        and(pr_and10[7],b[9],a[7]);


        and(pr_and10[8],b[9],a[8]);


        and(pr_and10[9],b[9],a[9]);


        and(pr_and10[10],b[9],a[10]);


        and(pr_and10[11],b[9],a[11]);


        and(pr_and10[12],b[9],a[12]);


        and(pr_and10[13],b[9],a[13]);


        and(pr_and10[14],b[9],a[14]);


        and(pr_and10[15],b[9],a[15]);


        and(pr_and10[16],b[9],a[16]);


        and(pr_and10[17],b[9],a[17]);


        and(pr_and10[18],b[9],a[18]);


        and(pr_and10[19],b[9],a[19]);


        and(pr_and10[20],b[9],a[20]);


        and(pr_and10[21],b[9],a[21]);


        and(pr_and10[22],b[9],a[22]);


        and(pr_and10[23],b[9],a[23]);


        and(pr_and10[24],b[9],a[24]);


        and(pr_and10[25],b[9],a[25]);


        and(pr_and10[26],b[9],a[26]);


        and(pr_and10[27],b[9],a[27]);


        and(pr_and10[28],b[9],a[28]);


        and(pr_and10[29],b[9],a[29]);


        and(pr_and10[30],b[9],a[30]);


        and(pr_and10[31],b[9],a[31]);


    not(si[9],pr_and10[31]);


        and(pr_and11[0],b[10],a[0]);


        and(pr_and11[1],b[10],a[1]);


        and(pr_and11[2],b[10],a[2]);


        and(pr_and11[3],b[10],a[3]);


        and(pr_and11[4],b[10],a[4]);


        and(pr_and11[5],b[10],a[5]);


        and(pr_and11[6],b[10],a[6]);


        and(pr_and11[7],b[10],a[7]);


        and(pr_and11[8],b[10],a[8]);


        and(pr_and11[9],b[10],a[9]);


        and(pr_and11[10],b[10],a[10]);


        and(pr_and11[11],b[10],a[11]);


        and(pr_and11[12],b[10],a[12]);


        and(pr_and11[13],b[10],a[13]);


        and(pr_and11[14],b[10],a[14]);


        and(pr_and11[15],b[10],a[15]);


        and(pr_and11[16],b[10],a[16]);


        and(pr_and11[17],b[10],a[17]);


        and(pr_and11[18],b[10],a[18]);


        and(pr_and11[19],b[10],a[19]);


        and(pr_and11[20],b[10],a[20]);


        and(pr_and11[21],b[10],a[21]);


        and(pr_and11[22],b[10],a[22]);


        and(pr_and11[23],b[10],a[23]);


        and(pr_and11[24],b[10],a[24]);


        and(pr_and11[25],b[10],a[25]);


        and(pr_and11[26],b[10],a[26]);


        and(pr_and11[27],b[10],a[27]);


        and(pr_and11[28],b[10],a[28]);


        and(pr_and11[29],b[10],a[29]);


        and(pr_and11[30],b[10],a[30]);


        and(pr_and11[31],b[10],a[31]);


    not(si[10],pr_and11[31]);


        and(pr_and12[0],b[11],a[0]);


        and(pr_and12[1],b[11],a[1]);


        and(pr_and12[2],b[11],a[2]);


        and(pr_and12[3],b[11],a[3]);


        and(pr_and12[4],b[11],a[4]);


        and(pr_and12[5],b[11],a[5]);


        and(pr_and12[6],b[11],a[6]);


        and(pr_and12[7],b[11],a[7]);


        and(pr_and12[8],b[11],a[8]);


        and(pr_and12[9],b[11],a[9]);


        and(pr_and12[10],b[11],a[10]);


        and(pr_and12[11],b[11],a[11]);


        and(pr_and12[12],b[11],a[12]);


        and(pr_and12[13],b[11],a[13]);


        and(pr_and12[14],b[11],a[14]);


        and(pr_and12[15],b[11],a[15]);


        and(pr_and12[16],b[11],a[16]);


        and(pr_and12[17],b[11],a[17]);


        and(pr_and12[18],b[11],a[18]);


        and(pr_and12[19],b[11],a[19]);


        and(pr_and12[20],b[11],a[20]);


        and(pr_and12[21],b[11],a[21]);


        and(pr_and12[22],b[11],a[22]);


        and(pr_and12[23],b[11],a[23]);


        and(pr_and12[24],b[11],a[24]);


        and(pr_and12[25],b[11],a[25]);


        and(pr_and12[26],b[11],a[26]);


        and(pr_and12[27],b[11],a[27]);


        and(pr_and12[28],b[11],a[28]);


        and(pr_and12[29],b[11],a[29]);


        and(pr_and12[30],b[11],a[30]);


        and(pr_and12[31],b[11],a[31]);


    not(si[11],pr_and12[31]);


        and(pr_and13[0],b[12],a[0]);


        and(pr_and13[1],b[12],a[1]);


        and(pr_and13[2],b[12],a[2]);


        and(pr_and13[3],b[12],a[3]);


        and(pr_and13[4],b[12],a[4]);


        and(pr_and13[5],b[12],a[5]);


        and(pr_and13[6],b[12],a[6]);


        and(pr_and13[7],b[12],a[7]);


        and(pr_and13[8],b[12],a[8]);


        and(pr_and13[9],b[12],a[9]);


        and(pr_and13[10],b[12],a[10]);


        and(pr_and13[11],b[12],a[11]);


        and(pr_and13[12],b[12],a[12]);


        and(pr_and13[13],b[12],a[13]);


        and(pr_and13[14],b[12],a[14]);


        and(pr_and13[15],b[12],a[15]);


        and(pr_and13[16],b[12],a[16]);


        and(pr_and13[17],b[12],a[17]);


        and(pr_and13[18],b[12],a[18]);


        and(pr_and13[19],b[12],a[19]);


        and(pr_and13[20],b[12],a[20]);


        and(pr_and13[21],b[12],a[21]);


        and(pr_and13[22],b[12],a[22]);


        and(pr_and13[23],b[12],a[23]);


        and(pr_and13[24],b[12],a[24]);


        and(pr_and13[25],b[12],a[25]);


        and(pr_and13[26],b[12],a[26]);


        and(pr_and13[27],b[12],a[27]);


        and(pr_and13[28],b[12],a[28]);


        and(pr_and13[29],b[12],a[29]);


        and(pr_and13[30],b[12],a[30]);


        and(pr_and13[31],b[12],a[31]);


    not(si[12],pr_and13[31]);


        and(pr_and14[0],b[13],a[0]);


        and(pr_and14[1],b[13],a[1]);


        and(pr_and14[2],b[13],a[2]);


        and(pr_and14[3],b[13],a[3]);


        and(pr_and14[4],b[13],a[4]);


        and(pr_and14[5],b[13],a[5]);


        and(pr_and14[6],b[13],a[6]);


        and(pr_and14[7],b[13],a[7]);


        and(pr_and14[8],b[13],a[8]);


        and(pr_and14[9],b[13],a[9]);


        and(pr_and14[10],b[13],a[10]);


        and(pr_and14[11],b[13],a[11]);


        and(pr_and14[12],b[13],a[12]);


        and(pr_and14[13],b[13],a[13]);


        and(pr_and14[14],b[13],a[14]);


        and(pr_and14[15],b[13],a[15]);


        and(pr_and14[16],b[13],a[16]);


        and(pr_and14[17],b[13],a[17]);


        and(pr_and14[18],b[13],a[18]);


        and(pr_and14[19],b[13],a[19]);


        and(pr_and14[20],b[13],a[20]);


        and(pr_and14[21],b[13],a[21]);


        and(pr_and14[22],b[13],a[22]);


        and(pr_and14[23],b[13],a[23]);


        and(pr_and14[24],b[13],a[24]);


        and(pr_and14[25],b[13],a[25]);


        and(pr_and14[26],b[13],a[26]);


        and(pr_and14[27],b[13],a[27]);


        and(pr_and14[28],b[13],a[28]);


        and(pr_and14[29],b[13],a[29]);


        and(pr_and14[30],b[13],a[30]);


        and(pr_and14[31],b[13],a[31]);


    not(si[13],pr_and14[31]);


        and(pr_and15[0],b[14],a[0]);


        and(pr_and15[1],b[14],a[1]);


        and(pr_and15[2],b[14],a[2]);


        and(pr_and15[3],b[14],a[3]);


        and(pr_and15[4],b[14],a[4]);


        and(pr_and15[5],b[14],a[5]);


        and(pr_and15[6],b[14],a[6]);


        and(pr_and15[7],b[14],a[7]);


        and(pr_and15[8],b[14],a[8]);


        and(pr_and15[9],b[14],a[9]);


        and(pr_and15[10],b[14],a[10]);


        and(pr_and15[11],b[14],a[11]);


        and(pr_and15[12],b[14],a[12]);


        and(pr_and15[13],b[14],a[13]);


        and(pr_and15[14],b[14],a[14]);


        and(pr_and15[15],b[14],a[15]);


        and(pr_and15[16],b[14],a[16]);


        and(pr_and15[17],b[14],a[17]);


        and(pr_and15[18],b[14],a[18]);


        and(pr_and15[19],b[14],a[19]);


        and(pr_and15[20],b[14],a[20]);


        and(pr_and15[21],b[14],a[21]);


        and(pr_and15[22],b[14],a[22]);


        and(pr_and15[23],b[14],a[23]);


        and(pr_and15[24],b[14],a[24]);


        and(pr_and15[25],b[14],a[25]);


        and(pr_and15[26],b[14],a[26]);


        and(pr_and15[27],b[14],a[27]);


        and(pr_and15[28],b[14],a[28]);


        and(pr_and15[29],b[14],a[29]);


        and(pr_and15[30],b[14],a[30]);


        and(pr_and15[31],b[14],a[31]);


    not(si[14],pr_and15[31]);


        and(pr_and16[0],b[15],a[0]);


        and(pr_and16[1],b[15],a[1]);


        and(pr_and16[2],b[15],a[2]);


        and(pr_and16[3],b[15],a[3]);


        and(pr_and16[4],b[15],a[4]);


        and(pr_and16[5],b[15],a[5]);


        and(pr_and16[6],b[15],a[6]);


        and(pr_and16[7],b[15],a[7]);


        and(pr_and16[8],b[15],a[8]);


        and(pr_and16[9],b[15],a[9]);


        and(pr_and16[10],b[15],a[10]);


        and(pr_and16[11],b[15],a[11]);


        and(pr_and16[12],b[15],a[12]);


        and(pr_and16[13],b[15],a[13]);


        and(pr_and16[14],b[15],a[14]);


        and(pr_and16[15],b[15],a[15]);


        and(pr_and16[16],b[15],a[16]);


        and(pr_and16[17],b[15],a[17]);


        and(pr_and16[18],b[15],a[18]);


        and(pr_and16[19],b[15],a[19]);


        and(pr_and16[20],b[15],a[20]);


        and(pr_and16[21],b[15],a[21]);


        and(pr_and16[22],b[15],a[22]);


        and(pr_and16[23],b[15],a[23]);


        and(pr_and16[24],b[15],a[24]);


        and(pr_and16[25],b[15],a[25]);


        and(pr_and16[26],b[15],a[26]);


        and(pr_and16[27],b[15],a[27]);


        and(pr_and16[28],b[15],a[28]);


        and(pr_and16[29],b[15],a[29]);


        and(pr_and16[30],b[15],a[30]);


        and(pr_and16[31],b[15],a[31]);


    not(si[15],pr_and16[31]);


        and(pr_and17[0],b[16],a[0]);


        and(pr_and17[1],b[16],a[1]);


        and(pr_and17[2],b[16],a[2]);


        and(pr_and17[3],b[16],a[3]);


        and(pr_and17[4],b[16],a[4]);


        and(pr_and17[5],b[16],a[5]);


        and(pr_and17[6],b[16],a[6]);


        and(pr_and17[7],b[16],a[7]);


        and(pr_and17[8],b[16],a[8]);


        and(pr_and17[9],b[16],a[9]);


        and(pr_and17[10],b[16],a[10]);


        and(pr_and17[11],b[16],a[11]);


        and(pr_and17[12],b[16],a[12]);


        and(pr_and17[13],b[16],a[13]);


        and(pr_and17[14],b[16],a[14]);


        and(pr_and17[15],b[16],a[15]);


        and(pr_and17[16],b[16],a[16]);


        and(pr_and17[17],b[16],a[17]);


        and(pr_and17[18],b[16],a[18]);


        and(pr_and17[19],b[16],a[19]);


        and(pr_and17[20],b[16],a[20]);


        and(pr_and17[21],b[16],a[21]);


        and(pr_and17[22],b[16],a[22]);


        and(pr_and17[23],b[16],a[23]);


        and(pr_and17[24],b[16],a[24]);


        and(pr_and17[25],b[16],a[25]);


        and(pr_and17[26],b[16],a[26]);


        and(pr_and17[27],b[16],a[27]);


        and(pr_and17[28],b[16],a[28]);


        and(pr_and17[29],b[16],a[29]);


        and(pr_and17[30],b[16],a[30]);


        and(pr_and17[31],b[16],a[31]);


    not(si[16],pr_and17[31]);


        and(pr_and18[0],b[17],a[0]);


        and(pr_and18[1],b[17],a[1]);


        and(pr_and18[2],b[17],a[2]);


        and(pr_and18[3],b[17],a[3]);


        and(pr_and18[4],b[17],a[4]);


        and(pr_and18[5],b[17],a[5]);


        and(pr_and18[6],b[17],a[6]);


        and(pr_and18[7],b[17],a[7]);


        and(pr_and18[8],b[17],a[8]);


        and(pr_and18[9],b[17],a[9]);


        and(pr_and18[10],b[17],a[10]);


        and(pr_and18[11],b[17],a[11]);


        and(pr_and18[12],b[17],a[12]);


        and(pr_and18[13],b[17],a[13]);


        and(pr_and18[14],b[17],a[14]);


        and(pr_and18[15],b[17],a[15]);


        and(pr_and18[16],b[17],a[16]);


        and(pr_and18[17],b[17],a[17]);


        and(pr_and18[18],b[17],a[18]);


        and(pr_and18[19],b[17],a[19]);


        and(pr_and18[20],b[17],a[20]);


        and(pr_and18[21],b[17],a[21]);


        and(pr_and18[22],b[17],a[22]);


        and(pr_and18[23],b[17],a[23]);


        and(pr_and18[24],b[17],a[24]);


        and(pr_and18[25],b[17],a[25]);


        and(pr_and18[26],b[17],a[26]);


        and(pr_and18[27],b[17],a[27]);


        and(pr_and18[28],b[17],a[28]);


        and(pr_and18[29],b[17],a[29]);


        and(pr_and18[30],b[17],a[30]);


        and(pr_and18[31],b[17],a[31]);


    not(si[17],pr_and18[31]);


        and(pr_and19[0],b[18],a[0]);


        and(pr_and19[1],b[18],a[1]);


        and(pr_and19[2],b[18],a[2]);


        and(pr_and19[3],b[18],a[3]);


        and(pr_and19[4],b[18],a[4]);


        and(pr_and19[5],b[18],a[5]);


        and(pr_and19[6],b[18],a[6]);


        and(pr_and19[7],b[18],a[7]);


        and(pr_and19[8],b[18],a[8]);


        and(pr_and19[9],b[18],a[9]);


        and(pr_and19[10],b[18],a[10]);


        and(pr_and19[11],b[18],a[11]);


        and(pr_and19[12],b[18],a[12]);


        and(pr_and19[13],b[18],a[13]);


        and(pr_and19[14],b[18],a[14]);


        and(pr_and19[15],b[18],a[15]);


        and(pr_and19[16],b[18],a[16]);


        and(pr_and19[17],b[18],a[17]);


        and(pr_and19[18],b[18],a[18]);


        and(pr_and19[19],b[18],a[19]);


        and(pr_and19[20],b[18],a[20]);


        and(pr_and19[21],b[18],a[21]);


        and(pr_and19[22],b[18],a[22]);


        and(pr_and19[23],b[18],a[23]);


        and(pr_and19[24],b[18],a[24]);


        and(pr_and19[25],b[18],a[25]);


        and(pr_and19[26],b[18],a[26]);


        and(pr_and19[27],b[18],a[27]);


        and(pr_and19[28],b[18],a[28]);


        and(pr_and19[29],b[18],a[29]);


        and(pr_and19[30],b[18],a[30]);


        and(pr_and19[31],b[18],a[31]);


    not(si[18],pr_and19[31]);


        and(pr_and20[0],b[19],a[0]);


        and(pr_and20[1],b[19],a[1]);


        and(pr_and20[2],b[19],a[2]);


        and(pr_and20[3],b[19],a[3]);


        and(pr_and20[4],b[19],a[4]);


        and(pr_and20[5],b[19],a[5]);


        and(pr_and20[6],b[19],a[6]);


        and(pr_and20[7],b[19],a[7]);


        and(pr_and20[8],b[19],a[8]);


        and(pr_and20[9],b[19],a[9]);


        and(pr_and20[10],b[19],a[10]);


        and(pr_and20[11],b[19],a[11]);


        and(pr_and20[12],b[19],a[12]);


        and(pr_and20[13],b[19],a[13]);


        and(pr_and20[14],b[19],a[14]);


        and(pr_and20[15],b[19],a[15]);


        and(pr_and20[16],b[19],a[16]);


        and(pr_and20[17],b[19],a[17]);


        and(pr_and20[18],b[19],a[18]);


        and(pr_and20[19],b[19],a[19]);


        and(pr_and20[20],b[19],a[20]);


        and(pr_and20[21],b[19],a[21]);


        and(pr_and20[22],b[19],a[22]);


        and(pr_and20[23],b[19],a[23]);


        and(pr_and20[24],b[19],a[24]);


        and(pr_and20[25],b[19],a[25]);


        and(pr_and20[26],b[19],a[26]);


        and(pr_and20[27],b[19],a[27]);


        and(pr_and20[28],b[19],a[28]);


        and(pr_and20[29],b[19],a[29]);


        and(pr_and20[30],b[19],a[30]);


        and(pr_and20[31],b[19],a[31]);


    not(si[19],pr_and20[31]);


        and(pr_and21[0],b[20],a[0]);


        and(pr_and21[1],b[20],a[1]);


        and(pr_and21[2],b[20],a[2]);


        and(pr_and21[3],b[20],a[3]);


        and(pr_and21[4],b[20],a[4]);


        and(pr_and21[5],b[20],a[5]);


        and(pr_and21[6],b[20],a[6]);


        and(pr_and21[7],b[20],a[7]);


        and(pr_and21[8],b[20],a[8]);


        and(pr_and21[9],b[20],a[9]);


        and(pr_and21[10],b[20],a[10]);


        and(pr_and21[11],b[20],a[11]);


        and(pr_and21[12],b[20],a[12]);


        and(pr_and21[13],b[20],a[13]);


        and(pr_and21[14],b[20],a[14]);


        and(pr_and21[15],b[20],a[15]);


        and(pr_and21[16],b[20],a[16]);


        and(pr_and21[17],b[20],a[17]);


        and(pr_and21[18],b[20],a[18]);


        and(pr_and21[19],b[20],a[19]);


        and(pr_and21[20],b[20],a[20]);


        and(pr_and21[21],b[20],a[21]);


        and(pr_and21[22],b[20],a[22]);


        and(pr_and21[23],b[20],a[23]);


        and(pr_and21[24],b[20],a[24]);


        and(pr_and21[25],b[20],a[25]);


        and(pr_and21[26],b[20],a[26]);


        and(pr_and21[27],b[20],a[27]);


        and(pr_and21[28],b[20],a[28]);


        and(pr_and21[29],b[20],a[29]);


        and(pr_and21[30],b[20],a[30]);


        and(pr_and21[31],b[20],a[31]);


    not(si[20],pr_and21[31]);


        and(pr_and22[0],b[21],a[0]);


        and(pr_and22[1],b[21],a[1]);


        and(pr_and22[2],b[21],a[2]);


        and(pr_and22[3],b[21],a[3]);


        and(pr_and22[4],b[21],a[4]);


        and(pr_and22[5],b[21],a[5]);


        and(pr_and22[6],b[21],a[6]);


        and(pr_and22[7],b[21],a[7]);


        and(pr_and22[8],b[21],a[8]);


        and(pr_and22[9],b[21],a[9]);


        and(pr_and22[10],b[21],a[10]);


        and(pr_and22[11],b[21],a[11]);


        and(pr_and22[12],b[21],a[12]);


        and(pr_and22[13],b[21],a[13]);


        and(pr_and22[14],b[21],a[14]);


        and(pr_and22[15],b[21],a[15]);


        and(pr_and22[16],b[21],a[16]);


        and(pr_and22[17],b[21],a[17]);


        and(pr_and22[18],b[21],a[18]);


        and(pr_and22[19],b[21],a[19]);


        and(pr_and22[20],b[21],a[20]);


        and(pr_and22[21],b[21],a[21]);


        and(pr_and22[22],b[21],a[22]);


        and(pr_and22[23],b[21],a[23]);


        and(pr_and22[24],b[21],a[24]);


        and(pr_and22[25],b[21],a[25]);


        and(pr_and22[26],b[21],a[26]);


        and(pr_and22[27],b[21],a[27]);


        and(pr_and22[28],b[21],a[28]);


        and(pr_and22[29],b[21],a[29]);


        and(pr_and22[30],b[21],a[30]);


        and(pr_and22[31],b[21],a[31]);


    not(si[21],pr_and22[31]);


        and(pr_and23[0],b[22],a[0]);


        and(pr_and23[1],b[22],a[1]);


        and(pr_and23[2],b[22],a[2]);


        and(pr_and23[3],b[22],a[3]);


        and(pr_and23[4],b[22],a[4]);


        and(pr_and23[5],b[22],a[5]);


        and(pr_and23[6],b[22],a[6]);


        and(pr_and23[7],b[22],a[7]);


        and(pr_and23[8],b[22],a[8]);


        and(pr_and23[9],b[22],a[9]);


        and(pr_and23[10],b[22],a[10]);


        and(pr_and23[11],b[22],a[11]);


        and(pr_and23[12],b[22],a[12]);


        and(pr_and23[13],b[22],a[13]);


        and(pr_and23[14],b[22],a[14]);


        and(pr_and23[15],b[22],a[15]);


        and(pr_and23[16],b[22],a[16]);


        and(pr_and23[17],b[22],a[17]);


        and(pr_and23[18],b[22],a[18]);


        and(pr_and23[19],b[22],a[19]);


        and(pr_and23[20],b[22],a[20]);


        and(pr_and23[21],b[22],a[21]);


        and(pr_and23[22],b[22],a[22]);


        and(pr_and23[23],b[22],a[23]);


        and(pr_and23[24],b[22],a[24]);


        and(pr_and23[25],b[22],a[25]);


        and(pr_and23[26],b[22],a[26]);


        and(pr_and23[27],b[22],a[27]);


        and(pr_and23[28],b[22],a[28]);


        and(pr_and23[29],b[22],a[29]);


        and(pr_and23[30],b[22],a[30]);


        and(pr_and23[31],b[22],a[31]);


    not(si[22],pr_and23[31]);


        and(pr_and24[0],b[23],a[0]);


        and(pr_and24[1],b[23],a[1]);


        and(pr_and24[2],b[23],a[2]);


        and(pr_and24[3],b[23],a[3]);


        and(pr_and24[4],b[23],a[4]);


        and(pr_and24[5],b[23],a[5]);


        and(pr_and24[6],b[23],a[6]);


        and(pr_and24[7],b[23],a[7]);


        and(pr_and24[8],b[23],a[8]);


        and(pr_and24[9],b[23],a[9]);


        and(pr_and24[10],b[23],a[10]);


        and(pr_and24[11],b[23],a[11]);


        and(pr_and24[12],b[23],a[12]);


        and(pr_and24[13],b[23],a[13]);


        and(pr_and24[14],b[23],a[14]);


        and(pr_and24[15],b[23],a[15]);


        and(pr_and24[16],b[23],a[16]);


        and(pr_and24[17],b[23],a[17]);


        and(pr_and24[18],b[23],a[18]);


        and(pr_and24[19],b[23],a[19]);


        and(pr_and24[20],b[23],a[20]);


        and(pr_and24[21],b[23],a[21]);


        and(pr_and24[22],b[23],a[22]);


        and(pr_and24[23],b[23],a[23]);


        and(pr_and24[24],b[23],a[24]);


        and(pr_and24[25],b[23],a[25]);


        and(pr_and24[26],b[23],a[26]);


        and(pr_and24[27],b[23],a[27]);


        and(pr_and24[28],b[23],a[28]);


        and(pr_and24[29],b[23],a[29]);


        and(pr_and24[30],b[23],a[30]);


        and(pr_and24[31],b[23],a[31]);


    not(si[23],pr_and24[31]);


        and(pr_and25[0],b[24],a[0]);


        and(pr_and25[1],b[24],a[1]);


        and(pr_and25[2],b[24],a[2]);


        and(pr_and25[3],b[24],a[3]);


        and(pr_and25[4],b[24],a[4]);


        and(pr_and25[5],b[24],a[5]);


        and(pr_and25[6],b[24],a[6]);


        and(pr_and25[7],b[24],a[7]);


        and(pr_and25[8],b[24],a[8]);


        and(pr_and25[9],b[24],a[9]);


        and(pr_and25[10],b[24],a[10]);


        and(pr_and25[11],b[24],a[11]);


        and(pr_and25[12],b[24],a[12]);


        and(pr_and25[13],b[24],a[13]);


        and(pr_and25[14],b[24],a[14]);


        and(pr_and25[15],b[24],a[15]);


        and(pr_and25[16],b[24],a[16]);


        and(pr_and25[17],b[24],a[17]);


        and(pr_and25[18],b[24],a[18]);


        and(pr_and25[19],b[24],a[19]);


        and(pr_and25[20],b[24],a[20]);


        and(pr_and25[21],b[24],a[21]);


        and(pr_and25[22],b[24],a[22]);


        and(pr_and25[23],b[24],a[23]);


        and(pr_and25[24],b[24],a[24]);


        and(pr_and25[25],b[24],a[25]);


        and(pr_and25[26],b[24],a[26]);


        and(pr_and25[27],b[24],a[27]);


        and(pr_and25[28],b[24],a[28]);


        and(pr_and25[29],b[24],a[29]);


        and(pr_and25[30],b[24],a[30]);


        and(pr_and25[31],b[24],a[31]);


    not(si[24],pr_and25[31]);


        and(pr_and26[0],b[25],a[0]);


        and(pr_and26[1],b[25],a[1]);


        and(pr_and26[2],b[25],a[2]);


        and(pr_and26[3],b[25],a[3]);


        and(pr_and26[4],b[25],a[4]);


        and(pr_and26[5],b[25],a[5]);


        and(pr_and26[6],b[25],a[6]);


        and(pr_and26[7],b[25],a[7]);


        and(pr_and26[8],b[25],a[8]);


        and(pr_and26[9],b[25],a[9]);


        and(pr_and26[10],b[25],a[10]);


        and(pr_and26[11],b[25],a[11]);


        and(pr_and26[12],b[25],a[12]);


        and(pr_and26[13],b[25],a[13]);


        and(pr_and26[14],b[25],a[14]);


        and(pr_and26[15],b[25],a[15]);


        and(pr_and26[16],b[25],a[16]);


        and(pr_and26[17],b[25],a[17]);


        and(pr_and26[18],b[25],a[18]);


        and(pr_and26[19],b[25],a[19]);


        and(pr_and26[20],b[25],a[20]);


        and(pr_and26[21],b[25],a[21]);


        and(pr_and26[22],b[25],a[22]);


        and(pr_and26[23],b[25],a[23]);


        and(pr_and26[24],b[25],a[24]);


        and(pr_and26[25],b[25],a[25]);


        and(pr_and26[26],b[25],a[26]);


        and(pr_and26[27],b[25],a[27]);


        and(pr_and26[28],b[25],a[28]);


        and(pr_and26[29],b[25],a[29]);


        and(pr_and26[30],b[25],a[30]);


        and(pr_and26[31],b[25],a[31]);


    not(si[25],pr_and26[31]);


        and(pr_and27[0],b[26],a[0]);


        and(pr_and27[1],b[26],a[1]);


        and(pr_and27[2],b[26],a[2]);


        and(pr_and27[3],b[26],a[3]);


        and(pr_and27[4],b[26],a[4]);


        and(pr_and27[5],b[26],a[5]);


        and(pr_and27[6],b[26],a[6]);


        and(pr_and27[7],b[26],a[7]);


        and(pr_and27[8],b[26],a[8]);


        and(pr_and27[9],b[26],a[9]);


        and(pr_and27[10],b[26],a[10]);


        and(pr_and27[11],b[26],a[11]);


        and(pr_and27[12],b[26],a[12]);


        and(pr_and27[13],b[26],a[13]);


        and(pr_and27[14],b[26],a[14]);


        and(pr_and27[15],b[26],a[15]);


        and(pr_and27[16],b[26],a[16]);


        and(pr_and27[17],b[26],a[17]);


        and(pr_and27[18],b[26],a[18]);


        and(pr_and27[19],b[26],a[19]);


        and(pr_and27[20],b[26],a[20]);


        and(pr_and27[21],b[26],a[21]);


        and(pr_and27[22],b[26],a[22]);


        and(pr_and27[23],b[26],a[23]);


        and(pr_and27[24],b[26],a[24]);


        and(pr_and27[25],b[26],a[25]);


        and(pr_and27[26],b[26],a[26]);


        and(pr_and27[27],b[26],a[27]);


        and(pr_and27[28],b[26],a[28]);


        and(pr_and27[29],b[26],a[29]);


        and(pr_and27[30],b[26],a[30]);


        and(pr_and27[31],b[26],a[31]);


    not(si[26],pr_and27[31]);


        and(pr_and28[0],b[27],a[0]);


        and(pr_and28[1],b[27],a[1]);


        and(pr_and28[2],b[27],a[2]);


        and(pr_and28[3],b[27],a[3]);


        and(pr_and28[4],b[27],a[4]);


        and(pr_and28[5],b[27],a[5]);


        and(pr_and28[6],b[27],a[6]);


        and(pr_and28[7],b[27],a[7]);


        and(pr_and28[8],b[27],a[8]);


        and(pr_and28[9],b[27],a[9]);


        and(pr_and28[10],b[27],a[10]);


        and(pr_and28[11],b[27],a[11]);


        and(pr_and28[12],b[27],a[12]);


        and(pr_and28[13],b[27],a[13]);


        and(pr_and28[14],b[27],a[14]);


        and(pr_and28[15],b[27],a[15]);


        and(pr_and28[16],b[27],a[16]);


        and(pr_and28[17],b[27],a[17]);


        and(pr_and28[18],b[27],a[18]);


        and(pr_and28[19],b[27],a[19]);


        and(pr_and28[20],b[27],a[20]);


        and(pr_and28[21],b[27],a[21]);


        and(pr_and28[22],b[27],a[22]);


        and(pr_and28[23],b[27],a[23]);


        and(pr_and28[24],b[27],a[24]);


        and(pr_and28[25],b[27],a[25]);


        and(pr_and28[26],b[27],a[26]);


        and(pr_and28[27],b[27],a[27]);


        and(pr_and28[28],b[27],a[28]);


        and(pr_and28[29],b[27],a[29]);


        and(pr_and28[30],b[27],a[30]);


        and(pr_and28[31],b[27],a[31]);


    not(si[27],pr_and28[31]);


        and(pr_and29[0],b[28],a[0]);


        and(pr_and29[1],b[28],a[1]);


        and(pr_and29[2],b[28],a[2]);


        and(pr_and29[3],b[28],a[3]);


        and(pr_and29[4],b[28],a[4]);


        and(pr_and29[5],b[28],a[5]);


        and(pr_and29[6],b[28],a[6]);


        and(pr_and29[7],b[28],a[7]);


        and(pr_and29[8],b[28],a[8]);


        and(pr_and29[9],b[28],a[9]);


        and(pr_and29[10],b[28],a[10]);


        and(pr_and29[11],b[28],a[11]);


        and(pr_and29[12],b[28],a[12]);


        and(pr_and29[13],b[28],a[13]);


        and(pr_and29[14],b[28],a[14]);


        and(pr_and29[15],b[28],a[15]);


        and(pr_and29[16],b[28],a[16]);


        and(pr_and29[17],b[28],a[17]);


        and(pr_and29[18],b[28],a[18]);


        and(pr_and29[19],b[28],a[19]);


        and(pr_and29[20],b[28],a[20]);


        and(pr_and29[21],b[28],a[21]);


        and(pr_and29[22],b[28],a[22]);


        and(pr_and29[23],b[28],a[23]);


        and(pr_and29[24],b[28],a[24]);


        and(pr_and29[25],b[28],a[25]);


        and(pr_and29[26],b[28],a[26]);


        and(pr_and29[27],b[28],a[27]);


        and(pr_and29[28],b[28],a[28]);


        and(pr_and29[29],b[28],a[29]);


        and(pr_and29[30],b[28],a[30]);


        and(pr_and29[31],b[28],a[31]);


    not(si[28],pr_and29[31]);


        and(pr_and30[0],b[29],a[0]);


        and(pr_and30[1],b[29],a[1]);


        and(pr_and30[2],b[29],a[2]);


        and(pr_and30[3],b[29],a[3]);


        and(pr_and30[4],b[29],a[4]);


        and(pr_and30[5],b[29],a[5]);


        and(pr_and30[6],b[29],a[6]);


        and(pr_and30[7],b[29],a[7]);


        and(pr_and30[8],b[29],a[8]);


        and(pr_and30[9],b[29],a[9]);


        and(pr_and30[10],b[29],a[10]);


        and(pr_and30[11],b[29],a[11]);


        and(pr_and30[12],b[29],a[12]);


        and(pr_and30[13],b[29],a[13]);


        and(pr_and30[14],b[29],a[14]);


        and(pr_and30[15],b[29],a[15]);


        and(pr_and30[16],b[29],a[16]);


        and(pr_and30[17],b[29],a[17]);


        and(pr_and30[18],b[29],a[18]);


        and(pr_and30[19],b[29],a[19]);


        and(pr_and30[20],b[29],a[20]);


        and(pr_and30[21],b[29],a[21]);


        and(pr_and30[22],b[29],a[22]);


        and(pr_and30[23],b[29],a[23]);


        and(pr_and30[24],b[29],a[24]);


        and(pr_and30[25],b[29],a[25]);


        and(pr_and30[26],b[29],a[26]);


        and(pr_and30[27],b[29],a[27]);


        and(pr_and30[28],b[29],a[28]);


        and(pr_and30[29],b[29],a[29]);


        and(pr_and30[30],b[29],a[30]);


        and(pr_and30[31],b[29],a[31]);


    not(si[29],pr_and30[31]);


        and(pr_and31[0],b[30],a[0]);


        and(pr_and31[1],b[30],a[1]);


        and(pr_and31[2],b[30],a[2]);


        and(pr_and31[3],b[30],a[3]);


        and(pr_and31[4],b[30],a[4]);


        and(pr_and31[5],b[30],a[5]);


        and(pr_and31[6],b[30],a[6]);


        and(pr_and31[7],b[30],a[7]);


        and(pr_and31[8],b[30],a[8]);


        and(pr_and31[9],b[30],a[9]);


        and(pr_and31[10],b[30],a[10]);


        and(pr_and31[11],b[30],a[11]);


        and(pr_and31[12],b[30],a[12]);


        and(pr_and31[13],b[30],a[13]);


        and(pr_and31[14],b[30],a[14]);


        and(pr_and31[15],b[30],a[15]);


        and(pr_and31[16],b[30],a[16]);


        and(pr_and31[17],b[30],a[17]);


        and(pr_and31[18],b[30],a[18]);


        and(pr_and31[19],b[30],a[19]);


        and(pr_and31[20],b[30],a[20]);


        and(pr_and31[21],b[30],a[21]);


        and(pr_and31[22],b[30],a[22]);


        and(pr_and31[23],b[30],a[23]);


        and(pr_and31[24],b[30],a[24]);


        and(pr_and31[25],b[30],a[25]);


        and(pr_and31[26],b[30],a[26]);


        and(pr_and31[27],b[30],a[27]);


        and(pr_and31[28],b[30],a[28]);


        and(pr_and31[29],b[30],a[29]);


        and(pr_and31[30],b[30],a[30]);


        and(pr_and31[31],b[30],a[31]);


    not(si[30],pr_and31[31]);


    and(pr_and32[0],b[31],~a[0]);

    and(pr_and32[1],b[31],~a[1]);

    and(pr_and32[2],b[31],~a[2]);

    and(pr_and32[3],b[31],~a[3]);

    and(pr_and32[4],b[31],~a[4]);

    and(pr_and32[5],b[31],~a[5]);

    and(pr_and32[6],b[31],~a[6]);

    and(pr_and32[7],b[31],~a[7]);

    and(pr_and32[8],b[31],~a[8]);

    and(pr_and32[9],b[31],~a[9]);

    and(pr_and32[10],b[31],~a[10]);

    and(pr_and32[11],b[31],~a[11]);

    and(pr_and32[12],b[31],~a[12]);

    and(pr_and32[13],b[31],~a[13]);

    and(pr_and32[14],b[31],~a[14]);

    and(pr_and32[15],b[31],~a[15]);

    and(pr_and32[16],b[31],~a[16]);

    and(pr_and32[17],b[31],~a[17]);

    and(pr_and32[18],b[31],~a[18]);

    and(pr_and32[19],b[31],~a[19]);

    and(pr_and32[20],b[31],~a[20]);

    and(pr_and32[21],b[31],~a[21]);

    and(pr_and32[22],b[31],~a[22]);

    and(pr_and32[23],b[31],~a[23]);

    and(pr_and32[24],b[31],~a[24]);

    and(pr_and32[25],b[31],~a[25]);

    and(pr_and32[26],b[31],~a[26]);

    and(pr_and32[27],b[31],~a[27]);

    and(pr_and32[28],b[31],~a[28]);

    and(pr_and32[29],b[31],~a[29]);

    and(pr_and32[30],b[31],~a[30]);

    and(pr_and32[31],b[31],~a[31]);

not(si[31],pr_and32[31]);


adder_half ha1(pr_and1[1],pr_and2[0],c1[0],p[1]);


adder_full fa1_1(pr_and1[2],pr_and2[1],pr_and3[0],c1[1],s1[0]);


adder_full fa1_2(pr_and1[3],pr_and2[2],pr_and3[1],c1[2],s1[1]);


adder_full fa1_3(pr_and1[4],pr_and2[3],pr_and3[2],c1[3],s1[2]);


adder_full fa1_4(pr_and1[5],pr_and2[4],pr_and3[3],c1[4],s1[3]);


adder_full fa1_5(pr_and1[6],pr_and2[5],pr_and3[4],c1[5],s1[4]);


adder_full fa1_6(pr_and1[7],pr_and2[6],pr_and3[5],c1[6],s1[5]);


adder_full fa1_7(pr_and1[8],pr_and2[7],pr_and3[6],c1[7],s1[6]);


adder_full fa1_8(pr_and1[9],pr_and2[8],pr_and3[7],c1[8],s1[7]);


adder_full fa1_9(pr_and1[10],pr_and2[9],pr_and3[8],c1[9],s1[8]);


adder_full fa1_10(pr_and1[11],pr_and2[10],pr_and3[9],c1[10],s1[9]);


adder_full fa1_11(pr_and1[12],pr_and2[11],pr_and3[10],c1[11],s1[10]);


adder_full fa1_12(pr_and1[13],pr_and2[12],pr_and3[11],c1[12],s1[11]);


adder_full fa1_13(pr_and1[14],pr_and2[13],pr_and3[12],c1[13],s1[12]);


adder_full fa1_14(pr_and1[15],pr_and2[14],pr_and3[13],c1[14],s1[13]);


adder_full fa1_15(pr_and1[16],pr_and2[15],pr_and3[14],c1[15],s1[14]);


adder_full fa1_16(pr_and1[17],pr_and2[16],pr_and3[15],c1[16],s1[15]);


adder_full fa1_17(pr_and1[18],pr_and2[17],pr_and3[16],c1[17],s1[16]);


adder_full fa1_18(pr_and1[19],pr_and2[18],pr_and3[17],c1[18],s1[17]);


adder_full fa1_19(pr_and1[20],pr_and2[19],pr_and3[18],c1[19],s1[18]);


adder_full fa1_20(pr_and1[21],pr_and2[20],pr_and3[19],c1[20],s1[19]);


adder_full fa1_21(pr_and1[22],pr_and2[21],pr_and3[20],c1[21],s1[20]);


adder_full fa1_22(pr_and1[23],pr_and2[22],pr_and3[21],c1[22],s1[21]);


adder_full fa1_23(pr_and1[24],pr_and2[23],pr_and3[22],c1[23],s1[22]);


adder_full fa1_24(pr_and1[25],pr_and2[24],pr_and3[23],c1[24],s1[23]);


adder_full fa1_25(pr_and1[26],pr_and2[25],pr_and3[24],c1[25],s1[24]);


adder_full fa1_26(pr_and1[27],pr_and2[26],pr_and3[25],c1[26],s1[25]);


adder_full fa1_27(pr_and1[28],pr_and2[27],pr_and3[26],c1[27],s1[26]);


adder_full fa1_28(pr_and1[29],pr_and2[28],pr_and3[27],c1[28],s1[27]);


adder_full fa1_29(pr_and1[30],pr_and2[29],pr_and3[28],c1[29],s1[28]);


adder_full fa1_30(pr_and1[31],pr_and2[30],pr_and3[29],c1[30],s1[29]);



adder_full fa2_31(si[0],si[1],pr_and3[30],c1[31],s1[30]);



//layer 2
adder_half ha2(s1[0],c1[0],c2[0],p[2]);


adder_full fa2_0(s1[1],c1[1],pr_and4[0],c2[1],s2[0]);


adder_full fa2_1(s1[2],c1[2],pr_and4[1],c2[2],s2[1]);


adder_full fa2_2(s1[3],c1[3],pr_and4[2],c2[3],s2[2]);


adder_full fa2_3(s1[4],c1[4],pr_and4[3],c2[4],s2[3]);


adder_full fa2_4(s1[5],c1[5],pr_and4[4],c2[5],s2[4]);


adder_full fa2_5(s1[6],c1[6],pr_and4[5],c2[6],s2[5]);


adder_full fa2_6(s1[7],c1[7],pr_and4[6],c2[7],s2[6]);


adder_full fa2_7(s1[8],c1[8],pr_and4[7],c2[8],s2[7]);


adder_full fa2_8(s1[9],c1[9],pr_and4[8],c2[9],s2[8]);


adder_full fa2_9(s1[10],c1[10],pr_and4[9],c2[10],s2[9]);


adder_full fa2_10(s1[11],c1[11],pr_and4[10],c2[11],s2[10]);


adder_full fa2_11(s1[12],c1[12],pr_and4[11],c2[12],s2[11]);


adder_full fa2_12(s1[13],c1[13],pr_and4[12],c2[13],s2[12]);


adder_full fa2_13(s1[14],c1[14],pr_and4[13],c2[14],s2[13]);


adder_full fa2_14(s1[15],c1[15],pr_and4[14],c2[15],s2[14]);


adder_full fa2_15(s1[16],c1[16],pr_and4[15],c2[16],s2[15]);


adder_full fa2_16(s1[17],c1[17],pr_and4[16],c2[17],s2[16]);


adder_full fa2_17(s1[18],c1[18],pr_and4[17],c2[18],s2[17]);


adder_full fa2_18(s1[19],c1[19],pr_and4[18],c2[19],s2[18]);


adder_full fa2_19(s1[20],c1[20],pr_and4[19],c2[20],s2[19]);


adder_full fa2_20(s1[21],c1[21],pr_and4[20],c2[21],s2[20]);


adder_full fa2_21(s1[22],c1[22],pr_and4[21],c2[22],s2[21]);


adder_full fa2_22(s1[23],c1[23],pr_and4[22],c2[23],s2[22]);


adder_full fa2_23(s1[24],c1[24],pr_and4[23],c2[24],s2[23]);


adder_full fa2_24(s1[25],c1[25],pr_and4[24],c2[25],s2[24]);


adder_full fa2_25(s1[26],c1[26],pr_and4[25],c2[26],s2[25]);


adder_full fa2_26(s1[27],c1[27],pr_and4[26],c2[27],s2[26]);


adder_full fa2_27(s1[28],c1[28],pr_and4[27],c2[28],s2[27]);


adder_full fa2_28(s1[29],c1[29],pr_and4[28],c2[29],s2[28]);


adder_full fa2_29(s1[30],c1[30],pr_and4[29],c2[30],s2[29]);


adder_full fa2_30(si[2],c1[31],pr_and4[30],c2[31],s2[30]);



//layer 3
adder_half ha3(s2[0],c2[0],c3[0],p[3]);


adder_full fa3_0(s2[1],c2[1],pr_and5[0],c3[1],s3[0]);


adder_full fa3_1(s2[2],c2[2],pr_and5[1],c3[2],s3[1]);


adder_full fa3_2(s2[3],c2[3],pr_and5[2],c3[3],s3[2]);


adder_full fa3_3(s2[4],c2[4],pr_and5[3],c3[4],s3[3]);


adder_full fa3_4(s2[5],c2[5],pr_and5[4],c3[5],s3[4]);


adder_full fa3_5(s2[6],c2[6],pr_and5[5],c3[6],s3[5]);


adder_full fa3_6(s2[7],c2[7],pr_and5[6],c3[7],s3[6]);


adder_full fa3_7(s2[8],c2[8],pr_and5[7],c3[8],s3[7]);


adder_full fa3_8(s2[9],c2[9],pr_and5[8],c3[9],s3[8]);


adder_full fa3_9(s2[10],c2[10],pr_and5[9],c3[10],s3[9]);


adder_full fa3_10(s2[11],c2[11],pr_and5[10],c3[11],s3[10]);


adder_full fa3_11(s2[12],c2[12],pr_and5[11],c3[12],s3[11]);


adder_full fa3_12(s2[13],c2[13],pr_and5[12],c3[13],s3[12]);


adder_full fa3_13(s2[14],c2[14],pr_and5[13],c3[14],s3[13]);


adder_full fa3_14(s2[15],c2[15],pr_and5[14],c3[15],s3[14]);


adder_full fa3_15(s2[16],c2[16],pr_and5[15],c3[16],s3[15]);


adder_full fa3_16(s2[17],c2[17],pr_and5[16],c3[17],s3[16]);


adder_full fa3_17(s2[18],c2[18],pr_and5[17],c3[18],s3[17]);


adder_full fa3_18(s2[19],c2[19],pr_and5[18],c3[19],s3[18]);


adder_full fa3_19(s2[20],c2[20],pr_and5[19],c3[20],s3[19]);


adder_full fa3_20(s2[21],c2[21],pr_and5[20],c3[21],s3[20]);


adder_full fa3_21(s2[22],c2[22],pr_and5[21],c3[22],s3[21]);


adder_full fa3_22(s2[23],c2[23],pr_and5[22],c3[23],s3[22]);


adder_full fa3_23(s2[24],c2[24],pr_and5[23],c3[24],s3[23]);


adder_full fa3_24(s2[25],c2[25],pr_and5[24],c3[25],s3[24]);


adder_full fa3_25(s2[26],c2[26],pr_and5[25],c3[26],s3[25]);


adder_full fa3_26(s2[27],c2[27],pr_and5[26],c3[27],s3[26]);


adder_full fa3_27(s2[28],c2[28],pr_and5[27],c3[28],s3[27]);


adder_full fa3_28(s2[29],c2[29],pr_and5[28],c3[29],s3[28]);


adder_full fa3_29(s2[30],c2[30],pr_and5[29],c3[30],s3[29]);


adder_full fa3_30(si[3],c2[31],pr_and5[30],c3[31],s3[30]);



//layer 4
adder_half ha4(s3[0],c3[0],c4[0],p[4]);


adder_full fa4_0(s3[1],c3[1],pr_and6[0],c4[1],s4[0]);


adder_full fa4_1(s3[2],c3[2],pr_and6[1],c4[2],s4[1]);


adder_full fa4_2(s3[3],c3[3],pr_and6[2],c4[3],s4[2]);


adder_full fa4_3(s3[4],c3[4],pr_and6[3],c4[4],s4[3]);


adder_full fa4_4(s3[5],c3[5],pr_and6[4],c4[5],s4[4]);


adder_full fa4_5(s3[6],c3[6],pr_and6[5],c4[6],s4[5]);


adder_full fa4_6(s3[7],c3[7],pr_and6[6],c4[7],s4[6]);


adder_full fa4_7(s3[8],c3[8],pr_and6[7],c4[8],s4[7]);


adder_full fa4_8(s3[9],c3[9],pr_and6[8],c4[9],s4[8]);


adder_full fa4_9(s3[10],c3[10],pr_and6[9],c4[10],s4[9]);


adder_full fa4_10(s3[11],c3[11],pr_and6[10],c4[11],s4[10]);


adder_full fa4_11(s3[12],c3[12],pr_and6[11],c4[12],s4[11]);


adder_full fa4_12(s3[13],c3[13],pr_and6[12],c4[13],s4[12]);


adder_full fa4_13(s3[14],c3[14],pr_and6[13],c4[14],s4[13]);


adder_full fa4_14(s3[15],c3[15],pr_and6[14],c4[15],s4[14]);


adder_full fa4_15(s3[16],c3[16],pr_and6[15],c4[16],s4[15]);


adder_full fa4_16(s3[17],c3[17],pr_and6[16],c4[17],s4[16]);


adder_full fa4_17(s3[18],c3[18],pr_and6[17],c4[18],s4[17]);


adder_full fa4_18(s3[19],c3[19],pr_and6[18],c4[19],s4[18]);


adder_full fa4_19(s3[20],c3[20],pr_and6[19],c4[20],s4[19]);


adder_full fa4_20(s3[21],c3[21],pr_and6[20],c4[21],s4[20]);


adder_full fa4_21(s3[22],c3[22],pr_and6[21],c4[22],s4[21]);


adder_full fa4_22(s3[23],c3[23],pr_and6[22],c4[23],s4[22]);


adder_full fa4_23(s3[24],c3[24],pr_and6[23],c4[24],s4[23]);


adder_full fa4_24(s3[25],c3[25],pr_and6[24],c4[25],s4[24]);


adder_full fa4_25(s3[26],c3[26],pr_and6[25],c4[26],s4[25]);


adder_full fa4_26(s3[27],c3[27],pr_and6[26],c4[27],s4[26]);


adder_full fa4_27(s3[28],c3[28],pr_and6[27],c4[28],s4[27]);


adder_full fa4_28(s3[29],c3[29],pr_and6[28],c4[29],s4[28]);


adder_full fa4_29(s3[30],c3[30],pr_and6[29],c4[30],s4[29]);


adder_full fa4_30(si[4],c3[31],pr_and6[30],c4[31],s4[30]);



//layer 5
adder_half ha5(s4[0],c4[0],c5[0],p[5]);


adder_full fa5_0(s4[1],c4[1],pr_and7[0],c5[1],s5[0]);


adder_full fa5_1(s4[2],c4[2],pr_and7[1],c5[2],s5[1]);


adder_full fa5_2(s4[3],c4[3],pr_and7[2],c5[3],s5[2]);


adder_full fa5_3(s4[4],c4[4],pr_and7[3],c5[4],s5[3]);


adder_full fa5_4(s4[5],c4[5],pr_and7[4],c5[5],s5[4]);


adder_full fa5_5(s4[6],c4[6],pr_and7[5],c5[6],s5[5]);


adder_full fa5_6(s4[7],c4[7],pr_and7[6],c5[7],s5[6]);


adder_full fa5_7(s4[8],c4[8],pr_and7[7],c5[8],s5[7]);


adder_full fa5_8(s4[9],c4[9],pr_and7[8],c5[9],s5[8]);


adder_full fa5_9(s4[10],c4[10],pr_and7[9],c5[10],s5[9]);


adder_full fa5_10(s4[11],c4[11],pr_and7[10],c5[11],s5[10]);


adder_full fa5_11(s4[12],c4[12],pr_and7[11],c5[12],s5[11]);


adder_full fa5_12(s4[13],c4[13],pr_and7[12],c5[13],s5[12]);


adder_full fa5_13(s4[14],c4[14],pr_and7[13],c5[14],s5[13]);


adder_full fa5_14(s4[15],c4[15],pr_and7[14],c5[15],s5[14]);


adder_full fa5_15(s4[16],c4[16],pr_and7[15],c5[16],s5[15]);


adder_full fa5_16(s4[17],c4[17],pr_and7[16],c5[17],s5[16]);


adder_full fa5_17(s4[18],c4[18],pr_and7[17],c5[18],s5[17]);


adder_full fa5_18(s4[19],c4[19],pr_and7[18],c5[19],s5[18]);


adder_full fa5_19(s4[20],c4[20],pr_and7[19],c5[20],s5[19]);


adder_full fa5_20(s4[21],c4[21],pr_and7[20],c5[21],s5[20]);


adder_full fa5_21(s4[22],c4[22],pr_and7[21],c5[22],s5[21]);


adder_full fa5_22(s4[23],c4[23],pr_and7[22],c5[23],s5[22]);


adder_full fa5_23(s4[24],c4[24],pr_and7[23],c5[24],s5[23]);


adder_full fa5_24(s4[25],c4[25],pr_and7[24],c5[25],s5[24]);


adder_full fa5_25(s4[26],c4[26],pr_and7[25],c5[26],s5[25]);


adder_full fa5_26(s4[27],c4[27],pr_and7[26],c5[27],s5[26]);


adder_full fa5_27(s4[28],c4[28],pr_and7[27],c5[28],s5[27]);


adder_full fa5_28(s4[29],c4[29],pr_and7[28],c5[29],s5[28]);


adder_full fa5_29(s4[30],c4[30],pr_and7[29],c5[30],s5[29]);


adder_full fa5_30(si[5],c4[31],pr_and7[30],c5[31],s5[30]);



//layer 6
adder_half ha6(s5[0],c5[0],c6[0],p[6]);


adder_full fa6_0(s5[1],c5[1],pr_and8[0],c6[1],s6[0]);


adder_full fa6_1(s5[2],c5[2],pr_and8[1],c6[2],s6[1]);


adder_full fa6_2(s5[3],c5[3],pr_and8[2],c6[3],s6[2]);


adder_full fa6_3(s5[4],c5[4],pr_and8[3],c6[4],s6[3]);


adder_full fa6_4(s5[5],c5[5],pr_and8[4],c6[5],s6[4]);


adder_full fa6_5(s5[6],c5[6],pr_and8[5],c6[6],s6[5]);


adder_full fa6_6(s5[7],c5[7],pr_and8[6],c6[7],s6[6]);


adder_full fa6_7(s5[8],c5[8],pr_and8[7],c6[8],s6[7]);


adder_full fa6_8(s5[9],c5[9],pr_and8[8],c6[9],s6[8]);


adder_full fa6_9(s5[10],c5[10],pr_and8[9],c6[10],s6[9]);


adder_full fa6_10(s5[11],c5[11],pr_and8[10],c6[11],s6[10]);


adder_full fa6_11(s5[12],c5[12],pr_and8[11],c6[12],s6[11]);


adder_full fa6_12(s5[13],c5[13],pr_and8[12],c6[13],s6[12]);


adder_full fa6_13(s5[14],c5[14],pr_and8[13],c6[14],s6[13]);


adder_full fa6_14(s5[15],c5[15],pr_and8[14],c6[15],s6[14]);


adder_full fa6_15(s5[16],c5[16],pr_and8[15],c6[16],s6[15]);


adder_full fa6_16(s5[17],c5[17],pr_and8[16],c6[17],s6[16]);


adder_full fa6_17(s5[18],c5[18],pr_and8[17],c6[18],s6[17]);


adder_full fa6_18(s5[19],c5[19],pr_and8[18],c6[19],s6[18]);


adder_full fa6_19(s5[20],c5[20],pr_and8[19],c6[20],s6[19]);


adder_full fa6_20(s5[21],c5[21],pr_and8[20],c6[21],s6[20]);


adder_full fa6_21(s5[22],c5[22],pr_and8[21],c6[22],s6[21]);


adder_full fa6_22(s5[23],c5[23],pr_and8[22],c6[23],s6[22]);


adder_full fa6_23(s5[24],c5[24],pr_and8[23],c6[24],s6[23]);


adder_full fa6_24(s5[25],c5[25],pr_and8[24],c6[25],s6[24]);


adder_full fa6_25(s5[26],c5[26],pr_and8[25],c6[26],s6[25]);


adder_full fa6_26(s5[27],c5[27],pr_and8[26],c6[27],s6[26]);


adder_full fa6_27(s5[28],c5[28],pr_and8[27],c6[28],s6[27]);


adder_full fa6_28(s5[29],c5[29],pr_and8[28],c6[29],s6[28]);


adder_full fa6_29(s5[30],c5[30],pr_and8[29],c6[30],s6[29]);


adder_full fa6_30(si[6],c5[31],pr_and8[30],c6[31],s6[30]);



//layer 7
adder_half ha7(s6[0],c6[0],c7[0],p[7]);


adder_full fa7_0(s6[1],c6[1],pr_and9[0],c7[1],s7[0]);


adder_full fa7_1(s6[2],c6[2],pr_and9[1],c7[2],s7[1]);


adder_full fa7_2(s6[3],c6[3],pr_and9[2],c7[3],s7[2]);


adder_full fa7_3(s6[4],c6[4],pr_and9[3],c7[4],s7[3]);


adder_full fa7_4(s6[5],c6[5],pr_and9[4],c7[5],s7[4]);


adder_full fa7_5(s6[6],c6[6],pr_and9[5],c7[6],s7[5]);


adder_full fa7_6(s6[7],c6[7],pr_and9[6],c7[7],s7[6]);


adder_full fa7_7(s6[8],c6[8],pr_and9[7],c7[8],s7[7]);


adder_full fa7_8(s6[9],c6[9],pr_and9[8],c7[9],s7[8]);


adder_full fa7_9(s6[10],c6[10],pr_and9[9],c7[10],s7[9]);


adder_full fa7_10(s6[11],c6[11],pr_and9[10],c7[11],s7[10]);


adder_full fa7_11(s6[12],c6[12],pr_and9[11],c7[12],s7[11]);


adder_full fa7_12(s6[13],c6[13],pr_and9[12],c7[13],s7[12]);


adder_full fa7_13(s6[14],c6[14],pr_and9[13],c7[14],s7[13]);


adder_full fa7_14(s6[15],c6[15],pr_and9[14],c7[15],s7[14]);


adder_full fa7_15(s6[16],c6[16],pr_and9[15],c7[16],s7[15]);


adder_full fa7_16(s6[17],c6[17],pr_and9[16],c7[17],s7[16]);


adder_full fa7_17(s6[18],c6[18],pr_and9[17],c7[18],s7[17]);


adder_full fa7_18(s6[19],c6[19],pr_and9[18],c7[19],s7[18]);


adder_full fa7_19(s6[20],c6[20],pr_and9[19],c7[20],s7[19]);


adder_full fa7_20(s6[21],c6[21],pr_and9[20],c7[21],s7[20]);


adder_full fa7_21(s6[22],c6[22],pr_and9[21],c7[22],s7[21]);


adder_full fa7_22(s6[23],c6[23],pr_and9[22],c7[23],s7[22]);


adder_full fa7_23(s6[24],c6[24],pr_and9[23],c7[24],s7[23]);


adder_full fa7_24(s6[25],c6[25],pr_and9[24],c7[25],s7[24]);


adder_full fa7_25(s6[26],c6[26],pr_and9[25],c7[26],s7[25]);


adder_full fa7_26(s6[27],c6[27],pr_and9[26],c7[27],s7[26]);


adder_full fa7_27(s6[28],c6[28],pr_and9[27],c7[28],s7[27]);


adder_full fa7_28(s6[29],c6[29],pr_and9[28],c7[29],s7[28]);


adder_full fa7_29(s6[30],c6[30],pr_and9[29],c7[30],s7[29]);


adder_full fa7_30(si[7],c6[31],pr_and9[30],c7[31],s7[30]);



//layer 8
adder_half ha8(s7[0],c7[0],c8[0],p[8]);


adder_full fa8_0(s7[1],c7[1],pr_and10[0],c8[1],s8[0]);


adder_full fa8_1(s7[2],c7[2],pr_and10[1],c8[2],s8[1]);


adder_full fa8_2(s7[3],c7[3],pr_and10[2],c8[3],s8[2]);


adder_full fa8_3(s7[4],c7[4],pr_and10[3],c8[4],s8[3]);


adder_full fa8_4(s7[5],c7[5],pr_and10[4],c8[5],s8[4]);


adder_full fa8_5(s7[6],c7[6],pr_and10[5],c8[6],s8[5]);


adder_full fa8_6(s7[7],c7[7],pr_and10[6],c8[7],s8[6]);


adder_full fa8_7(s7[8],c7[8],pr_and10[7],c8[8],s8[7]);


adder_full fa8_8(s7[9],c7[9],pr_and10[8],c8[9],s8[8]);


adder_full fa8_9(s7[10],c7[10],pr_and10[9],c8[10],s8[9]);


adder_full fa8_10(s7[11],c7[11],pr_and10[10],c8[11],s8[10]);


adder_full fa8_11(s7[12],c7[12],pr_and10[11],c8[12],s8[11]);


adder_full fa8_12(s7[13],c7[13],pr_and10[12],c8[13],s8[12]);


adder_full fa8_13(s7[14],c7[14],pr_and10[13],c8[14],s8[13]);


adder_full fa8_14(s7[15],c7[15],pr_and10[14],c8[15],s8[14]);


adder_full fa8_15(s7[16],c7[16],pr_and10[15],c8[16],s8[15]);


adder_full fa8_16(s7[17],c7[17],pr_and10[16],c8[17],s8[16]);


adder_full fa8_17(s7[18],c7[18],pr_and10[17],c8[18],s8[17]);


adder_full fa8_18(s7[19],c7[19],pr_and10[18],c8[19],s8[18]);


adder_full fa8_19(s7[20],c7[20],pr_and10[19],c8[20],s8[19]);


adder_full fa8_20(s7[21],c7[21],pr_and10[20],c8[21],s8[20]);


adder_full fa8_21(s7[22],c7[22],pr_and10[21],c8[22],s8[21]);


adder_full fa8_22(s7[23],c7[23],pr_and10[22],c8[23],s8[22]);


adder_full fa8_23(s7[24],c7[24],pr_and10[23],c8[24],s8[23]);


adder_full fa8_24(s7[25],c7[25],pr_and10[24],c8[25],s8[24]);


adder_full fa8_25(s7[26],c7[26],pr_and10[25],c8[26],s8[25]);


adder_full fa8_26(s7[27],c7[27],pr_and10[26],c8[27],s8[26]);


adder_full fa8_27(s7[28],c7[28],pr_and10[27],c8[28],s8[27]);


adder_full fa8_28(s7[29],c7[29],pr_and10[28],c8[29],s8[28]);


adder_full fa8_29(s7[30],c7[30],pr_and10[29],c8[30],s8[29]);


adder_full fa8_30(si[8],c7[31],pr_and10[30],c8[31],s8[30]);



//layer 9
adder_half ha9(s8[0],c8[0],c9[0],p[9]);


adder_full fa9_0(s8[1],c8[1],pr_and11[0],c9[1],s9[0]);


adder_full fa9_1(s8[2],c8[2],pr_and11[1],c9[2],s9[1]);


adder_full fa9_2(s8[3],c8[3],pr_and11[2],c9[3],s9[2]);


adder_full fa9_3(s8[4],c8[4],pr_and11[3],c9[4],s9[3]);


adder_full fa9_4(s8[5],c8[5],pr_and11[4],c9[5],s9[4]);


adder_full fa9_5(s8[6],c8[6],pr_and11[5],c9[6],s9[5]);


adder_full fa9_6(s8[7],c8[7],pr_and11[6],c9[7],s9[6]);


adder_full fa9_7(s8[8],c8[8],pr_and11[7],c9[8],s9[7]);


adder_full fa9_8(s8[9],c8[9],pr_and11[8],c9[9],s9[8]);


adder_full fa9_9(s8[10],c8[10],pr_and11[9],c9[10],s9[9]);


adder_full fa9_10(s8[11],c8[11],pr_and11[10],c9[11],s9[10]);


adder_full fa9_11(s8[12],c8[12],pr_and11[11],c9[12],s9[11]);


adder_full fa9_12(s8[13],c8[13],pr_and11[12],c9[13],s9[12]);


adder_full fa9_13(s8[14],c8[14],pr_and11[13],c9[14],s9[13]);


adder_full fa9_14(s8[15],c8[15],pr_and11[14],c9[15],s9[14]);


adder_full fa9_15(s8[16],c8[16],pr_and11[15],c9[16],s9[15]);


adder_full fa9_16(s8[17],c8[17],pr_and11[16],c9[17],s9[16]);


adder_full fa9_17(s8[18],c8[18],pr_and11[17],c9[18],s9[17]);


adder_full fa9_18(s8[19],c8[19],pr_and11[18],c9[19],s9[18]);


adder_full fa9_19(s8[20],c8[20],pr_and11[19],c9[20],s9[19]);


adder_full fa9_20(s8[21],c8[21],pr_and11[20],c9[21],s9[20]);


adder_full fa9_21(s8[22],c8[22],pr_and11[21],c9[22],s9[21]);


adder_full fa9_22(s8[23],c8[23],pr_and11[22],c9[23],s9[22]);


adder_full fa9_23(s8[24],c8[24],pr_and11[23],c9[24],s9[23]);


adder_full fa9_24(s8[25],c8[25],pr_and11[24],c9[25],s9[24]);


adder_full fa9_25(s8[26],c8[26],pr_and11[25],c9[26],s9[25]);


adder_full fa9_26(s8[27],c8[27],pr_and11[26],c9[27],s9[26]);


adder_full fa9_27(s8[28],c8[28],pr_and11[27],c9[28],s9[27]);


adder_full fa9_28(s8[29],c8[29],pr_and11[28],c9[29],s9[28]);


adder_full fa9_29(s8[30],c8[30],pr_and11[29],c9[30],s9[29]);


adder_full fa9_30(si[9],c8[31],pr_and11[30],c9[31],s9[30]);



//layer 10
adder_half ha10(s9[0],c9[0],c10[0],p[10]);


adder_full fa10_0(s9[1],c9[1],pr_and12[0],c10[1],s10[0]);


adder_full fa10_1(s9[2],c9[2],pr_and12[1],c10[2],s10[1]);


adder_full fa10_2(s9[3],c9[3],pr_and12[2],c10[3],s10[2]);


adder_full fa10_3(s9[4],c9[4],pr_and12[3],c10[4],s10[3]);


adder_full fa10_4(s9[5],c9[5],pr_and12[4],c10[5],s10[4]);


adder_full fa10_5(s9[6],c9[6],pr_and12[5],c10[6],s10[5]);


adder_full fa10_6(s9[7],c9[7],pr_and12[6],c10[7],s10[6]);


adder_full fa10_7(s9[8],c9[8],pr_and12[7],c10[8],s10[7]);


adder_full fa10_8(s9[9],c9[9],pr_and12[8],c10[9],s10[8]);


adder_full fa10_9(s9[10],c9[10],pr_and12[9],c10[10],s10[9]);


adder_full fa10_10(s9[11],c9[11],pr_and12[10],c10[11],s10[10]);


adder_full fa10_11(s9[12],c9[12],pr_and12[11],c10[12],s10[11]);


adder_full fa10_12(s9[13],c9[13],pr_and12[12],c10[13],s10[12]);


adder_full fa10_13(s9[14],c9[14],pr_and12[13],c10[14],s10[13]);


adder_full fa10_14(s9[15],c9[15],pr_and12[14],c10[15],s10[14]);


adder_full fa10_15(s9[16],c9[16],pr_and12[15],c10[16],s10[15]);


adder_full fa10_16(s9[17],c9[17],pr_and12[16],c10[17],s10[16]);


adder_full fa10_17(s9[18],c9[18],pr_and12[17],c10[18],s10[17]);


adder_full fa10_18(s9[19],c9[19],pr_and12[18],c10[19],s10[18]);


adder_full fa10_19(s9[20],c9[20],pr_and12[19],c10[20],s10[19]);


adder_full fa10_20(s9[21],c9[21],pr_and12[20],c10[21],s10[20]);


adder_full fa10_21(s9[22],c9[22],pr_and12[21],c10[22],s10[21]);


adder_full fa10_22(s9[23],c9[23],pr_and12[22],c10[23],s10[22]);


adder_full fa10_23(s9[24],c9[24],pr_and12[23],c10[24],s10[23]);


adder_full fa10_24(s9[25],c9[25],pr_and12[24],c10[25],s10[24]);


adder_full fa10_25(s9[26],c9[26],pr_and12[25],c10[26],s10[25]);


adder_full fa10_26(s9[27],c9[27],pr_and12[26],c10[27],s10[26]);


adder_full fa10_27(s9[28],c9[28],pr_and12[27],c10[28],s10[27]);


adder_full fa10_28(s9[29],c9[29],pr_and12[28],c10[29],s10[28]);


adder_full fa10_29(s9[30],c9[30],pr_and12[29],c10[30],s10[29]);


adder_full fa10_30(si[10],c9[31],pr_and12[30],c10[31],s10[30]);



//layer 11
adder_half ha11(s10[0],c10[0],c11[0],p[11]);


adder_full fa11_0(s10[1],c10[1],pr_and13[0],c11[1],s11[0]);


adder_full fa11_1(s10[2],c10[2],pr_and13[1],c11[2],s11[1]);


adder_full fa11_2(s10[3],c10[3],pr_and13[2],c11[3],s11[2]);


adder_full fa11_3(s10[4],c10[4],pr_and13[3],c11[4],s11[3]);


adder_full fa11_4(s10[5],c10[5],pr_and13[4],c11[5],s11[4]);


adder_full fa11_5(s10[6],c10[6],pr_and13[5],c11[6],s11[5]);


adder_full fa11_6(s10[7],c10[7],pr_and13[6],c11[7],s11[6]);


adder_full fa11_7(s10[8],c10[8],pr_and13[7],c11[8],s11[7]);


adder_full fa11_8(s10[9],c10[9],pr_and13[8],c11[9],s11[8]);


adder_full fa11_9(s10[10],c10[10],pr_and13[9],c11[10],s11[9]);


adder_full fa11_10(s10[11],c10[11],pr_and13[10],c11[11],s11[10]);


adder_full fa11_11(s10[12],c10[12],pr_and13[11],c11[12],s11[11]);


adder_full fa11_12(s10[13],c10[13],pr_and13[12],c11[13],s11[12]);


adder_full fa11_13(s10[14],c10[14],pr_and13[13],c11[14],s11[13]);


adder_full fa11_14(s10[15],c10[15],pr_and13[14],c11[15],s11[14]);


adder_full fa11_15(s10[16],c10[16],pr_and13[15],c11[16],s11[15]);


adder_full fa11_16(s10[17],c10[17],pr_and13[16],c11[17],s11[16]);


adder_full fa11_17(s10[18],c10[18],pr_and13[17],c11[18],s11[17]);


adder_full fa11_18(s10[19],c10[19],pr_and13[18],c11[19],s11[18]);


adder_full fa11_19(s10[20],c10[20],pr_and13[19],c11[20],s11[19]);


adder_full fa11_20(s10[21],c10[21],pr_and13[20],c11[21],s11[20]);


adder_full fa11_21(s10[22],c10[22],pr_and13[21],c11[22],s11[21]);


adder_full fa11_22(s10[23],c10[23],pr_and13[22],c11[23],s11[22]);


adder_full fa11_23(s10[24],c10[24],pr_and13[23],c11[24],s11[23]);


adder_full fa11_24(s10[25],c10[25],pr_and13[24],c11[25],s11[24]);


adder_full fa11_25(s10[26],c10[26],pr_and13[25],c11[26],s11[25]);


adder_full fa11_26(s10[27],c10[27],pr_and13[26],c11[27],s11[26]);


adder_full fa11_27(s10[28],c10[28],pr_and13[27],c11[28],s11[27]);


adder_full fa11_28(s10[29],c10[29],pr_and13[28],c11[29],s11[28]);


adder_full fa11_29(s10[30],c10[30],pr_and13[29],c11[30],s11[29]);


adder_full fa11_30(si[11],c10[31],pr_and13[30],c11[31],s11[30]);



//layer 12
adder_half ha12(s11[0],c11[0],c12[0],p[12]);


adder_full fa12_0(s11[1],c11[1],pr_and14[0],c12[1],s12[0]);


adder_full fa12_1(s11[2],c11[2],pr_and14[1],c12[2],s12[1]);


adder_full fa12_2(s11[3],c11[3],pr_and14[2],c12[3],s12[2]);


adder_full fa12_3(s11[4],c11[4],pr_and14[3],c12[4],s12[3]);


adder_full fa12_4(s11[5],c11[5],pr_and14[4],c12[5],s12[4]);


adder_full fa12_5(s11[6],c11[6],pr_and14[5],c12[6],s12[5]);


adder_full fa12_6(s11[7],c11[7],pr_and14[6],c12[7],s12[6]);


adder_full fa12_7(s11[8],c11[8],pr_and14[7],c12[8],s12[7]);


adder_full fa12_8(s11[9],c11[9],pr_and14[8],c12[9],s12[8]);


adder_full fa12_9(s11[10],c11[10],pr_and14[9],c12[10],s12[9]);


adder_full fa12_10(s11[11],c11[11],pr_and14[10],c12[11],s12[10]);


adder_full fa12_11(s11[12],c11[12],pr_and14[11],c12[12],s12[11]);


adder_full fa12_12(s11[13],c11[13],pr_and14[12],c12[13],s12[12]);


adder_full fa12_13(s11[14],c11[14],pr_and14[13],c12[14],s12[13]);


adder_full fa12_14(s11[15],c11[15],pr_and14[14],c12[15],s12[14]);


adder_full fa12_15(s11[16],c11[16],pr_and14[15],c12[16],s12[15]);


adder_full fa12_16(s11[17],c11[17],pr_and14[16],c12[17],s12[16]);


adder_full fa12_17(s11[18],c11[18],pr_and14[17],c12[18],s12[17]);


adder_full fa12_18(s11[19],c11[19],pr_and14[18],c12[19],s12[18]);


adder_full fa12_19(s11[20],c11[20],pr_and14[19],c12[20],s12[19]);


adder_full fa12_20(s11[21],c11[21],pr_and14[20],c12[21],s12[20]);


adder_full fa12_21(s11[22],c11[22],pr_and14[21],c12[22],s12[21]);


adder_full fa12_22(s11[23],c11[23],pr_and14[22],c12[23],s12[22]);


adder_full fa12_23(s11[24],c11[24],pr_and14[23],c12[24],s12[23]);


adder_full fa12_24(s11[25],c11[25],pr_and14[24],c12[25],s12[24]);


adder_full fa12_25(s11[26],c11[26],pr_and14[25],c12[26],s12[25]);


adder_full fa12_26(s11[27],c11[27],pr_and14[26],c12[27],s12[26]);


adder_full fa12_27(s11[28],c11[28],pr_and14[27],c12[28],s12[27]);


adder_full fa12_28(s11[29],c11[29],pr_and14[28],c12[29],s12[28]);


adder_full fa12_29(s11[30],c11[30],pr_and14[29],c12[30],s12[29]);


adder_full fa12_30(si[12],c11[31],pr_and14[30],c12[31],s12[30]);



//layer 13
adder_half ha13(s12[0],c12[0],c13[0],p[13]);


adder_full fa13_0(s12[1],c12[1],pr_and15[0],c13[1],s13[0]);


adder_full fa13_1(s12[2],c12[2],pr_and15[1],c13[2],s13[1]);


adder_full fa13_2(s12[3],c12[3],pr_and15[2],c13[3],s13[2]);


adder_full fa13_3(s12[4],c12[4],pr_and15[3],c13[4],s13[3]);


adder_full fa13_4(s12[5],c12[5],pr_and15[4],c13[5],s13[4]);


adder_full fa13_5(s12[6],c12[6],pr_and15[5],c13[6],s13[5]);


adder_full fa13_6(s12[7],c12[7],pr_and15[6],c13[7],s13[6]);


adder_full fa13_7(s12[8],c12[8],pr_and15[7],c13[8],s13[7]);


adder_full fa13_8(s12[9],c12[9],pr_and15[8],c13[9],s13[8]);


adder_full fa13_9(s12[10],c12[10],pr_and15[9],c13[10],s13[9]);


adder_full fa13_10(s12[11],c12[11],pr_and15[10],c13[11],s13[10]);


adder_full fa13_11(s12[12],c12[12],pr_and15[11],c13[12],s13[11]);


adder_full fa13_12(s12[13],c12[13],pr_and15[12],c13[13],s13[12]);


adder_full fa13_13(s12[14],c12[14],pr_and15[13],c13[14],s13[13]);


adder_full fa13_14(s12[15],c12[15],pr_and15[14],c13[15],s13[14]);


adder_full fa13_15(s12[16],c12[16],pr_and15[15],c13[16],s13[15]);


adder_full fa13_16(s12[17],c12[17],pr_and15[16],c13[17],s13[16]);


adder_full fa13_17(s12[18],c12[18],pr_and15[17],c13[18],s13[17]);


adder_full fa13_18(s12[19],c12[19],pr_and15[18],c13[19],s13[18]);


adder_full fa13_19(s12[20],c12[20],pr_and15[19],c13[20],s13[19]);


adder_full fa13_20(s12[21],c12[21],pr_and15[20],c13[21],s13[20]);


adder_full fa13_21(s12[22],c12[22],pr_and15[21],c13[22],s13[21]);


adder_full fa13_22(s12[23],c12[23],pr_and15[22],c13[23],s13[22]);


adder_full fa13_23(s12[24],c12[24],pr_and15[23],c13[24],s13[23]);


adder_full fa13_24(s12[25],c12[25],pr_and15[24],c13[25],s13[24]);


adder_full fa13_25(s12[26],c12[26],pr_and15[25],c13[26],s13[25]);


adder_full fa13_26(s12[27],c12[27],pr_and15[26],c13[27],s13[26]);


adder_full fa13_27(s12[28],c12[28],pr_and15[27],c13[28],s13[27]);


adder_full fa13_28(s12[29],c12[29],pr_and15[28],c13[29],s13[28]);


adder_full fa13_29(s12[30],c12[30],pr_and15[29],c13[30],s13[29]);


adder_full fa13_30(si[13],c12[31],pr_and15[30],c13[31],s13[30]);



//layer 14
adder_half ha14(s13[0],c13[0],c14[0],p[14]);


adder_full fa14_0(s13[1],c13[1],pr_and16[0],c14[1],s14[0]);


adder_full fa14_1(s13[2],c13[2],pr_and16[1],c14[2],s14[1]);


adder_full fa14_2(s13[3],c13[3],pr_and16[2],c14[3],s14[2]);


adder_full fa14_3(s13[4],c13[4],pr_and16[3],c14[4],s14[3]);


adder_full fa14_4(s13[5],c13[5],pr_and16[4],c14[5],s14[4]);


adder_full fa14_5(s13[6],c13[6],pr_and16[5],c14[6],s14[5]);


adder_full fa14_6(s13[7],c13[7],pr_and16[6],c14[7],s14[6]);


adder_full fa14_7(s13[8],c13[8],pr_and16[7],c14[8],s14[7]);


adder_full fa14_8(s13[9],c13[9],pr_and16[8],c14[9],s14[8]);


adder_full fa14_9(s13[10],c13[10],pr_and16[9],c14[10],s14[9]);


adder_full fa14_10(s13[11],c13[11],pr_and16[10],c14[11],s14[10]);


adder_full fa14_11(s13[12],c13[12],pr_and16[11],c14[12],s14[11]);


adder_full fa14_12(s13[13],c13[13],pr_and16[12],c14[13],s14[12]);


adder_full fa14_13(s13[14],c13[14],pr_and16[13],c14[14],s14[13]);


adder_full fa14_14(s13[15],c13[15],pr_and16[14],c14[15],s14[14]);


adder_full fa14_15(s13[16],c13[16],pr_and16[15],c14[16],s14[15]);


adder_full fa14_16(s13[17],c13[17],pr_and16[16],c14[17],s14[16]);


adder_full fa14_17(s13[18],c13[18],pr_and16[17],c14[18],s14[17]);


adder_full fa14_18(s13[19],c13[19],pr_and16[18],c14[19],s14[18]);


adder_full fa14_19(s13[20],c13[20],pr_and16[19],c14[20],s14[19]);


adder_full fa14_20(s13[21],c13[21],pr_and16[20],c14[21],s14[20]);


adder_full fa14_21(s13[22],c13[22],pr_and16[21],c14[22],s14[21]);


adder_full fa14_22(s13[23],c13[23],pr_and16[22],c14[23],s14[22]);


adder_full fa14_23(s13[24],c13[24],pr_and16[23],c14[24],s14[23]);


adder_full fa14_24(s13[25],c13[25],pr_and16[24],c14[25],s14[24]);


adder_full fa14_25(s13[26],c13[26],pr_and16[25],c14[26],s14[25]);


adder_full fa14_26(s13[27],c13[27],pr_and16[26],c14[27],s14[26]);


adder_full fa14_27(s13[28],c13[28],pr_and16[27],c14[28],s14[27]);


adder_full fa14_28(s13[29],c13[29],pr_and16[28],c14[29],s14[28]);


adder_full fa14_29(s13[30],c13[30],pr_and16[29],c14[30],s14[29]);


adder_full fa14_30(si[14],c13[31],pr_and16[30],c14[31],s14[30]);



//layer 15
adder_half ha15(s14[0],c14[0],c15[0],p[15]);


adder_full fa15_0(s14[1],c14[1],pr_and17[0],c15[1],s15[0]);


adder_full fa15_1(s14[2],c14[2],pr_and17[1],c15[2],s15[1]);


adder_full fa15_2(s14[3],c14[3],pr_and17[2],c15[3],s15[2]);


adder_full fa15_3(s14[4],c14[4],pr_and17[3],c15[4],s15[3]);


adder_full fa15_4(s14[5],c14[5],pr_and17[4],c15[5],s15[4]);


adder_full fa15_5(s14[6],c14[6],pr_and17[5],c15[6],s15[5]);


adder_full fa15_6(s14[7],c14[7],pr_and17[6],c15[7],s15[6]);


adder_full fa15_7(s14[8],c14[8],pr_and17[7],c15[8],s15[7]);


adder_full fa15_8(s14[9],c14[9],pr_and17[8],c15[9],s15[8]);


adder_full fa15_9(s14[10],c14[10],pr_and17[9],c15[10],s15[9]);


adder_full fa15_10(s14[11],c14[11],pr_and17[10],c15[11],s15[10]);


adder_full fa15_11(s14[12],c14[12],pr_and17[11],c15[12],s15[11]);


adder_full fa15_12(s14[13],c14[13],pr_and17[12],c15[13],s15[12]);


adder_full fa15_13(s14[14],c14[14],pr_and17[13],c15[14],s15[13]);


adder_full fa15_14(s14[15],c14[15],pr_and17[14],c15[15],s15[14]);


adder_full fa15_15(s14[16],c14[16],pr_and17[15],c15[16],s15[15]);


adder_full fa15_16(s14[17],c14[17],pr_and17[16],c15[17],s15[16]);


adder_full fa15_17(s14[18],c14[18],pr_and17[17],c15[18],s15[17]);


adder_full fa15_18(s14[19],c14[19],pr_and17[18],c15[19],s15[18]);


adder_full fa15_19(s14[20],c14[20],pr_and17[19],c15[20],s15[19]);


adder_full fa15_20(s14[21],c14[21],pr_and17[20],c15[21],s15[20]);


adder_full fa15_21(s14[22],c14[22],pr_and17[21],c15[22],s15[21]);


adder_full fa15_22(s14[23],c14[23],pr_and17[22],c15[23],s15[22]);


adder_full fa15_23(s14[24],c14[24],pr_and17[23],c15[24],s15[23]);


adder_full fa15_24(s14[25],c14[25],pr_and17[24],c15[25],s15[24]);


adder_full fa15_25(s14[26],c14[26],pr_and17[25],c15[26],s15[25]);


adder_full fa15_26(s14[27],c14[27],pr_and17[26],c15[27],s15[26]);


adder_full fa15_27(s14[28],c14[28],pr_and17[27],c15[28],s15[27]);


adder_full fa15_28(s14[29],c14[29],pr_and17[28],c15[29],s15[28]);


adder_full fa15_29(s14[30],c14[30],pr_and17[29],c15[30],s15[29]);


adder_full fa15_30(si[15],c14[31],pr_and17[30],c15[31],s15[30]);



//layer 16
adder_half ha16(s15[0],c15[0],c16[0],p[16]);


adder_full fa16_0(s15[1],c15[1],pr_and18[0],c16[1],s16[0]);


adder_full fa16_1(s15[2],c15[2],pr_and18[1],c16[2],s16[1]);


adder_full fa16_2(s15[3],c15[3],pr_and18[2],c16[3],s16[2]);


adder_full fa16_3(s15[4],c15[4],pr_and18[3],c16[4],s16[3]);


adder_full fa16_4(s15[5],c15[5],pr_and18[4],c16[5],s16[4]);


adder_full fa16_5(s15[6],c15[6],pr_and18[5],c16[6],s16[5]);


adder_full fa16_6(s15[7],c15[7],pr_and18[6],c16[7],s16[6]);


adder_full fa16_7(s15[8],c15[8],pr_and18[7],c16[8],s16[7]);


adder_full fa16_8(s15[9],c15[9],pr_and18[8],c16[9],s16[8]);


adder_full fa16_9(s15[10],c15[10],pr_and18[9],c16[10],s16[9]);


adder_full fa16_10(s15[11],c15[11],pr_and18[10],c16[11],s16[10]);


adder_full fa16_11(s15[12],c15[12],pr_and18[11],c16[12],s16[11]);


adder_full fa16_12(s15[13],c15[13],pr_and18[12],c16[13],s16[12]);


adder_full fa16_13(s15[14],c15[14],pr_and18[13],c16[14],s16[13]);


adder_full fa16_14(s15[15],c15[15],pr_and18[14],c16[15],s16[14]);


adder_full fa16_15(s15[16],c15[16],pr_and18[15],c16[16],s16[15]);


adder_full fa16_16(s15[17],c15[17],pr_and18[16],c16[17],s16[16]);


adder_full fa16_17(s15[18],c15[18],pr_and18[17],c16[18],s16[17]);


adder_full fa16_18(s15[19],c15[19],pr_and18[18],c16[19],s16[18]);


adder_full fa16_19(s15[20],c15[20],pr_and18[19],c16[20],s16[19]);


adder_full fa16_20(s15[21],c15[21],pr_and18[20],c16[21],s16[20]);


adder_full fa16_21(s15[22],c15[22],pr_and18[21],c16[22],s16[21]);


adder_full fa16_22(s15[23],c15[23],pr_and18[22],c16[23],s16[22]);


adder_full fa16_23(s15[24],c15[24],pr_and18[23],c16[24],s16[23]);


adder_full fa16_24(s15[25],c15[25],pr_and18[24],c16[25],s16[24]);


adder_full fa16_25(s15[26],c15[26],pr_and18[25],c16[26],s16[25]);


adder_full fa16_26(s15[27],c15[27],pr_and18[26],c16[27],s16[26]);


adder_full fa16_27(s15[28],c15[28],pr_and18[27],c16[28],s16[27]);


adder_full fa16_28(s15[29],c15[29],pr_and18[28],c16[29],s16[28]);


adder_full fa16_29(s15[30],c15[30],pr_and18[29],c16[30],s16[29]);


adder_full fa16_30(si[16],c15[31],pr_and18[30],c16[31],s16[30]);



//layer 17
adder_half ha17(s16[0],c16[0],c17[0],p[17]);


adder_full fa17_0(s16[1],c16[1],pr_and19[0],c17[1],s17[0]);


adder_full fa17_1(s16[2],c16[2],pr_and19[1],c17[2],s17[1]);


adder_full fa17_2(s16[3],c16[3],pr_and19[2],c17[3],s17[2]);


adder_full fa17_3(s16[4],c16[4],pr_and19[3],c17[4],s17[3]);


adder_full fa17_4(s16[5],c16[5],pr_and19[4],c17[5],s17[4]);


adder_full fa17_5(s16[6],c16[6],pr_and19[5],c17[6],s17[5]);


adder_full fa17_6(s16[7],c16[7],pr_and19[6],c17[7],s17[6]);


adder_full fa17_7(s16[8],c16[8],pr_and19[7],c17[8],s17[7]);


adder_full fa17_8(s16[9],c16[9],pr_and19[8],c17[9],s17[8]);


adder_full fa17_9(s16[10],c16[10],pr_and19[9],c17[10],s17[9]);


adder_full fa17_10(s16[11],c16[11],pr_and19[10],c17[11],s17[10]);


adder_full fa17_11(s16[12],c16[12],pr_and19[11],c17[12],s17[11]);


adder_full fa17_12(s16[13],c16[13],pr_and19[12],c17[13],s17[12]);


adder_full fa17_13(s16[14],c16[14],pr_and19[13],c17[14],s17[13]);


adder_full fa17_14(s16[15],c16[15],pr_and19[14],c17[15],s17[14]);


adder_full fa17_15(s16[16],c16[16],pr_and19[15],c17[16],s17[15]);


adder_full fa17_16(s16[17],c16[17],pr_and19[16],c17[17],s17[16]);


adder_full fa17_17(s16[18],c16[18],pr_and19[17],c17[18],s17[17]);


adder_full fa17_18(s16[19],c16[19],pr_and19[18],c17[19],s17[18]);


adder_full fa17_19(s16[20],c16[20],pr_and19[19],c17[20],s17[19]);


adder_full fa17_20(s16[21],c16[21],pr_and19[20],c17[21],s17[20]);


adder_full fa17_21(s16[22],c16[22],pr_and19[21],c17[22],s17[21]);


adder_full fa17_22(s16[23],c16[23],pr_and19[22],c17[23],s17[22]);


adder_full fa17_23(s16[24],c16[24],pr_and19[23],c17[24],s17[23]);


adder_full fa17_24(s16[25],c16[25],pr_and19[24],c17[25],s17[24]);


adder_full fa17_25(s16[26],c16[26],pr_and19[25],c17[26],s17[25]);


adder_full fa17_26(s16[27],c16[27],pr_and19[26],c17[27],s17[26]);


adder_full fa17_27(s16[28],c16[28],pr_and19[27],c17[28],s17[27]);


adder_full fa17_28(s16[29],c16[29],pr_and19[28],c17[29],s17[28]);


adder_full fa17_29(s16[30],c16[30],pr_and19[29],c17[30],s17[29]);


adder_full fa17_30(si[17],c16[31],pr_and19[30],c17[31],s17[30]);



//layer 18
adder_half ha18(s17[0],c17[0],c18[0],p[18]);


adder_full fa18_0(s17[1],c17[1],pr_and20[0],c18[1],s18[0]);


adder_full fa18_1(s17[2],c17[2],pr_and20[1],c18[2],s18[1]);


adder_full fa18_2(s17[3],c17[3],pr_and20[2],c18[3],s18[2]);


adder_full fa18_3(s17[4],c17[4],pr_and20[3],c18[4],s18[3]);


adder_full fa18_4(s17[5],c17[5],pr_and20[4],c18[5],s18[4]);


adder_full fa18_5(s17[6],c17[6],pr_and20[5],c18[6],s18[5]);


adder_full fa18_6(s17[7],c17[7],pr_and20[6],c18[7],s18[6]);


adder_full fa18_7(s17[8],c17[8],pr_and20[7],c18[8],s18[7]);


adder_full fa18_8(s17[9],c17[9],pr_and20[8],c18[9],s18[8]);


adder_full fa18_9(s17[10],c17[10],pr_and20[9],c18[10],s18[9]);


adder_full fa18_10(s17[11],c17[11],pr_and20[10],c18[11],s18[10]);


adder_full fa18_11(s17[12],c17[12],pr_and20[11],c18[12],s18[11]);


adder_full fa18_12(s17[13],c17[13],pr_and20[12],c18[13],s18[12]);


adder_full fa18_13(s17[14],c17[14],pr_and20[13],c18[14],s18[13]);


adder_full fa18_14(s17[15],c17[15],pr_and20[14],c18[15],s18[14]);


adder_full fa18_15(s17[16],c17[16],pr_and20[15],c18[16],s18[15]);


adder_full fa18_16(s17[17],c17[17],pr_and20[16],c18[17],s18[16]);


adder_full fa18_17(s17[18],c17[18],pr_and20[17],c18[18],s18[17]);


adder_full fa18_18(s17[19],c17[19],pr_and20[18],c18[19],s18[18]);


adder_full fa18_19(s17[20],c17[20],pr_and20[19],c18[20],s18[19]);


adder_full fa18_20(s17[21],c17[21],pr_and20[20],c18[21],s18[20]);


adder_full fa18_21(s17[22],c17[22],pr_and20[21],c18[22],s18[21]);


adder_full fa18_22(s17[23],c17[23],pr_and20[22],c18[23],s18[22]);


adder_full fa18_23(s17[24],c17[24],pr_and20[23],c18[24],s18[23]);


adder_full fa18_24(s17[25],c17[25],pr_and20[24],c18[25],s18[24]);


adder_full fa18_25(s17[26],c17[26],pr_and20[25],c18[26],s18[25]);


adder_full fa18_26(s17[27],c17[27],pr_and20[26],c18[27],s18[26]);


adder_full fa18_27(s17[28],c17[28],pr_and20[27],c18[28],s18[27]);


adder_full fa18_28(s17[29],c17[29],pr_and20[28],c18[29],s18[28]);


adder_full fa18_29(s17[30],c17[30],pr_and20[29],c18[30],s18[29]);


adder_full fa18_30(si[18],c17[31],pr_and20[30],c18[31],s18[30]);



//layer 19
adder_half ha19(s18[0],c18[0],c19[0],p[19]);


adder_full fa19_0(s18[1],c18[1],pr_and21[0],c19[1],s19[0]);


adder_full fa19_1(s18[2],c18[2],pr_and21[1],c19[2],s19[1]);


adder_full fa19_2(s18[3],c18[3],pr_and21[2],c19[3],s19[2]);


adder_full fa19_3(s18[4],c18[4],pr_and21[3],c19[4],s19[3]);


adder_full fa19_4(s18[5],c18[5],pr_and21[4],c19[5],s19[4]);


adder_full fa19_5(s18[6],c18[6],pr_and21[5],c19[6],s19[5]);


adder_full fa19_6(s18[7],c18[7],pr_and21[6],c19[7],s19[6]);


adder_full fa19_7(s18[8],c18[8],pr_and21[7],c19[8],s19[7]);


adder_full fa19_8(s18[9],c18[9],pr_and21[8],c19[9],s19[8]);


adder_full fa19_9(s18[10],c18[10],pr_and21[9],c19[10],s19[9]);


adder_full fa19_10(s18[11],c18[11],pr_and21[10],c19[11],s19[10]);


adder_full fa19_11(s18[12],c18[12],pr_and21[11],c19[12],s19[11]);


adder_full fa19_12(s18[13],c18[13],pr_and21[12],c19[13],s19[12]);


adder_full fa19_13(s18[14],c18[14],pr_and21[13],c19[14],s19[13]);


adder_full fa19_14(s18[15],c18[15],pr_and21[14],c19[15],s19[14]);


adder_full fa19_15(s18[16],c18[16],pr_and21[15],c19[16],s19[15]);


adder_full fa19_16(s18[17],c18[17],pr_and21[16],c19[17],s19[16]);


adder_full fa19_17(s18[18],c18[18],pr_and21[17],c19[18],s19[17]);


adder_full fa19_18(s18[19],c18[19],pr_and21[18],c19[19],s19[18]);


adder_full fa19_19(s18[20],c18[20],pr_and21[19],c19[20],s19[19]);


adder_full fa19_20(s18[21],c18[21],pr_and21[20],c19[21],s19[20]);


adder_full fa19_21(s18[22],c18[22],pr_and21[21],c19[22],s19[21]);


adder_full fa19_22(s18[23],c18[23],pr_and21[22],c19[23],s19[22]);


adder_full fa19_23(s18[24],c18[24],pr_and21[23],c19[24],s19[23]);


adder_full fa19_24(s18[25],c18[25],pr_and21[24],c19[25],s19[24]);


adder_full fa19_25(s18[26],c18[26],pr_and21[25],c19[26],s19[25]);


adder_full fa19_26(s18[27],c18[27],pr_and21[26],c19[27],s19[26]);


adder_full fa19_27(s18[28],c18[28],pr_and21[27],c19[28],s19[27]);


adder_full fa19_28(s18[29],c18[29],pr_and21[28],c19[29],s19[28]);


adder_full fa19_29(s18[30],c18[30],pr_and21[29],c19[30],s19[29]);


adder_full fa19_30(si[19],c18[31],pr_and21[30],c19[31],s19[30]);



//layer 20
adder_half ha20(s19[0],c19[0],c20[0],p[20]);


adder_full fa20_0(s19[1],c19[1],pr_and22[0],c20[1],s20[0]);


adder_full fa20_1(s19[2],c19[2],pr_and22[1],c20[2],s20[1]);


adder_full fa20_2(s19[3],c19[3],pr_and22[2],c20[3],s20[2]);


adder_full fa20_3(s19[4],c19[4],pr_and22[3],c20[4],s20[3]);


adder_full fa20_4(s19[5],c19[5],pr_and22[4],c20[5],s20[4]);


adder_full fa20_5(s19[6],c19[6],pr_and22[5],c20[6],s20[5]);


adder_full fa20_6(s19[7],c19[7],pr_and22[6],c20[7],s20[6]);


adder_full fa20_7(s19[8],c19[8],pr_and22[7],c20[8],s20[7]);


adder_full fa20_8(s19[9],c19[9],pr_and22[8],c20[9],s20[8]);


adder_full fa20_9(s19[10],c19[10],pr_and22[9],c20[10],s20[9]);


adder_full fa20_10(s19[11],c19[11],pr_and22[10],c20[11],s20[10]);


adder_full fa20_11(s19[12],c19[12],pr_and22[11],c20[12],s20[11]);


adder_full fa20_12(s19[13],c19[13],pr_and22[12],c20[13],s20[12]);


adder_full fa20_13(s19[14],c19[14],pr_and22[13],c20[14],s20[13]);


adder_full fa20_14(s19[15],c19[15],pr_and22[14],c20[15],s20[14]);


adder_full fa20_15(s19[16],c19[16],pr_and22[15],c20[16],s20[15]);


adder_full fa20_16(s19[17],c19[17],pr_and22[16],c20[17],s20[16]);


adder_full fa20_17(s19[18],c19[18],pr_and22[17],c20[18],s20[17]);


adder_full fa20_18(s19[19],c19[19],pr_and22[18],c20[19],s20[18]);


adder_full fa20_19(s19[20],c19[20],pr_and22[19],c20[20],s20[19]);


adder_full fa20_20(s19[21],c19[21],pr_and22[20],c20[21],s20[20]);


adder_full fa20_21(s19[22],c19[22],pr_and22[21],c20[22],s20[21]);


adder_full fa20_22(s19[23],c19[23],pr_and22[22],c20[23],s20[22]);


adder_full fa20_23(s19[24],c19[24],pr_and22[23],c20[24],s20[23]);


adder_full fa20_24(s19[25],c19[25],pr_and22[24],c20[25],s20[24]);


adder_full fa20_25(s19[26],c19[26],pr_and22[25],c20[26],s20[25]);


adder_full fa20_26(s19[27],c19[27],pr_and22[26],c20[27],s20[26]);


adder_full fa20_27(s19[28],c19[28],pr_and22[27],c20[28],s20[27]);


adder_full fa20_28(s19[29],c19[29],pr_and22[28],c20[29],s20[28]);


adder_full fa20_29(s19[30],c19[30],pr_and22[29],c20[30],s20[29]);


adder_full fa20_30(si[20],c19[31],pr_and22[30],c20[31],s20[30]);



//layer 21
adder_half ha21(s20[0],c20[0],c21[0],p[21]);


adder_full fa21_0(s20[1],c20[1],pr_and23[0],c21[1],s21[0]);


adder_full fa21_1(s20[2],c20[2],pr_and23[1],c21[2],s21[1]);


adder_full fa21_2(s20[3],c20[3],pr_and23[2],c21[3],s21[2]);


adder_full fa21_3(s20[4],c20[4],pr_and23[3],c21[4],s21[3]);


adder_full fa21_4(s20[5],c20[5],pr_and23[4],c21[5],s21[4]);


adder_full fa21_5(s20[6],c20[6],pr_and23[5],c21[6],s21[5]);


adder_full fa21_6(s20[7],c20[7],pr_and23[6],c21[7],s21[6]);


adder_full fa21_7(s20[8],c20[8],pr_and23[7],c21[8],s21[7]);


adder_full fa21_8(s20[9],c20[9],pr_and23[8],c21[9],s21[8]);


adder_full fa21_9(s20[10],c20[10],pr_and23[9],c21[10],s21[9]);


adder_full fa21_10(s20[11],c20[11],pr_and23[10],c21[11],s21[10]);


adder_full fa21_11(s20[12],c20[12],pr_and23[11],c21[12],s21[11]);


adder_full fa21_12(s20[13],c20[13],pr_and23[12],c21[13],s21[12]);


adder_full fa21_13(s20[14],c20[14],pr_and23[13],c21[14],s21[13]);


adder_full fa21_14(s20[15],c20[15],pr_and23[14],c21[15],s21[14]);


adder_full fa21_15(s20[16],c20[16],pr_and23[15],c21[16],s21[15]);


adder_full fa21_16(s20[17],c20[17],pr_and23[16],c21[17],s21[16]);


adder_full fa21_17(s20[18],c20[18],pr_and23[17],c21[18],s21[17]);


adder_full fa21_18(s20[19],c20[19],pr_and23[18],c21[19],s21[18]);


adder_full fa21_19(s20[20],c20[20],pr_and23[19],c21[20],s21[19]);


adder_full fa21_20(s20[21],c20[21],pr_and23[20],c21[21],s21[20]);


adder_full fa21_21(s20[22],c20[22],pr_and23[21],c21[22],s21[21]);


adder_full fa21_22(s20[23],c20[23],pr_and23[22],c21[23],s21[22]);


adder_full fa21_23(s20[24],c20[24],pr_and23[23],c21[24],s21[23]);


adder_full fa21_24(s20[25],c20[25],pr_and23[24],c21[25],s21[24]);


adder_full fa21_25(s20[26],c20[26],pr_and23[25],c21[26],s21[25]);


adder_full fa21_26(s20[27],c20[27],pr_and23[26],c21[27],s21[26]);


adder_full fa21_27(s20[28],c20[28],pr_and23[27],c21[28],s21[27]);


adder_full fa21_28(s20[29],c20[29],pr_and23[28],c21[29],s21[28]);


adder_full fa21_29(s20[30],c20[30],pr_and23[29],c21[30],s21[29]);


adder_full fa21_30(si[21],c20[31],pr_and23[30],c21[31],s21[30]);



//layer 22
adder_half ha22(s21[0],c21[0],c22[0],p[22]);


adder_full fa22_0(s21[1],c21[1],pr_and24[0],c22[1],s22[0]);


adder_full fa22_1(s21[2],c21[2],pr_and24[1],c22[2],s22[1]);


adder_full fa22_2(s21[3],c21[3],pr_and24[2],c22[3],s22[2]);


adder_full fa22_3(s21[4],c21[4],pr_and24[3],c22[4],s22[3]);


adder_full fa22_4(s21[5],c21[5],pr_and24[4],c22[5],s22[4]);


adder_full fa22_5(s21[6],c21[6],pr_and24[5],c22[6],s22[5]);


adder_full fa22_6(s21[7],c21[7],pr_and24[6],c22[7],s22[6]);


adder_full fa22_7(s21[8],c21[8],pr_and24[7],c22[8],s22[7]);


adder_full fa22_8(s21[9],c21[9],pr_and24[8],c22[9],s22[8]);


adder_full fa22_9(s21[10],c21[10],pr_and24[9],c22[10],s22[9]);


adder_full fa22_10(s21[11],c21[11],pr_and24[10],c22[11],s22[10]);


adder_full fa22_11(s21[12],c21[12],pr_and24[11],c22[12],s22[11]);


adder_full fa22_12(s21[13],c21[13],pr_and24[12],c22[13],s22[12]);


adder_full fa22_13(s21[14],c21[14],pr_and24[13],c22[14],s22[13]);


adder_full fa22_14(s21[15],c21[15],pr_and24[14],c22[15],s22[14]);


adder_full fa22_15(s21[16],c21[16],pr_and24[15],c22[16],s22[15]);


adder_full fa22_16(s21[17],c21[17],pr_and24[16],c22[17],s22[16]);


adder_full fa22_17(s21[18],c21[18],pr_and24[17],c22[18],s22[17]);


adder_full fa22_18(s21[19],c21[19],pr_and24[18],c22[19],s22[18]);


adder_full fa22_19(s21[20],c21[20],pr_and24[19],c22[20],s22[19]);


adder_full fa22_20(s21[21],c21[21],pr_and24[20],c22[21],s22[20]);


adder_full fa22_21(s21[22],c21[22],pr_and24[21],c22[22],s22[21]);


adder_full fa22_22(s21[23],c21[23],pr_and24[22],c22[23],s22[22]);


adder_full fa22_23(s21[24],c21[24],pr_and24[23],c22[24],s22[23]);


adder_full fa22_24(s21[25],c21[25],pr_and24[24],c22[25],s22[24]);


adder_full fa22_25(s21[26],c21[26],pr_and24[25],c22[26],s22[25]);


adder_full fa22_26(s21[27],c21[27],pr_and24[26],c22[27],s22[26]);


adder_full fa22_27(s21[28],c21[28],pr_and24[27],c22[28],s22[27]);


adder_full fa22_28(s21[29],c21[29],pr_and24[28],c22[29],s22[28]);


adder_full fa22_29(s21[30],c21[30],pr_and24[29],c22[30],s22[29]);


adder_full fa22_30(si[22],c21[31],pr_and24[30],c22[31],s22[30]);



//layer 23
adder_half ha23(s22[0],c22[0],c23[0],p[23]);


adder_full fa23_0(s22[1],c22[1],pr_and25[0],c23[1],s23[0]);


adder_full fa23_1(s22[2],c22[2],pr_and25[1],c23[2],s23[1]);


adder_full fa23_2(s22[3],c22[3],pr_and25[2],c23[3],s23[2]);


adder_full fa23_3(s22[4],c22[4],pr_and25[3],c23[4],s23[3]);


adder_full fa23_4(s22[5],c22[5],pr_and25[4],c23[5],s23[4]);


adder_full fa23_5(s22[6],c22[6],pr_and25[5],c23[6],s23[5]);


adder_full fa23_6(s22[7],c22[7],pr_and25[6],c23[7],s23[6]);


adder_full fa23_7(s22[8],c22[8],pr_and25[7],c23[8],s23[7]);


adder_full fa23_8(s22[9],c22[9],pr_and25[8],c23[9],s23[8]);


adder_full fa23_9(s22[10],c22[10],pr_and25[9],c23[10],s23[9]);


adder_full fa23_10(s22[11],c22[11],pr_and25[10],c23[11],s23[10]);


adder_full fa23_11(s22[12],c22[12],pr_and25[11],c23[12],s23[11]);


adder_full fa23_12(s22[13],c22[13],pr_and25[12],c23[13],s23[12]);


adder_full fa23_13(s22[14],c22[14],pr_and25[13],c23[14],s23[13]);


adder_full fa23_14(s22[15],c22[15],pr_and25[14],c23[15],s23[14]);


adder_full fa23_15(s22[16],c22[16],pr_and25[15],c23[16],s23[15]);


adder_full fa23_16(s22[17],c22[17],pr_and25[16],c23[17],s23[16]);


adder_full fa23_17(s22[18],c22[18],pr_and25[17],c23[18],s23[17]);


adder_full fa23_18(s22[19],c22[19],pr_and25[18],c23[19],s23[18]);


adder_full fa23_19(s22[20],c22[20],pr_and25[19],c23[20],s23[19]);


adder_full fa23_20(s22[21],c22[21],pr_and25[20],c23[21],s23[20]);


adder_full fa23_21(s22[22],c22[22],pr_and25[21],c23[22],s23[21]);


adder_full fa23_22(s22[23],c22[23],pr_and25[22],c23[23],s23[22]);


adder_full fa23_23(s22[24],c22[24],pr_and25[23],c23[24],s23[23]);


adder_full fa23_24(s22[25],c22[25],pr_and25[24],c23[25],s23[24]);


adder_full fa23_25(s22[26],c22[26],pr_and25[25],c23[26],s23[25]);


adder_full fa23_26(s22[27],c22[27],pr_and25[26],c23[27],s23[26]);


adder_full fa23_27(s22[28],c22[28],pr_and25[27],c23[28],s23[27]);


adder_full fa23_28(s22[29],c22[29],pr_and25[28],c23[29],s23[28]);


adder_full fa23_29(s22[30],c22[30],pr_and25[29],c23[30],s23[29]);


adder_full fa23_30(si[23],c22[31],pr_and25[30],c23[31],s23[30]);



//layer 24
adder_half ha24(s23[0],c23[0],c24[0],p[24]);


adder_full fa24_0(s23[1],c23[1],pr_and26[0],c24[1],s24[0]);


adder_full fa24_1(s23[2],c23[2],pr_and26[1],c24[2],s24[1]);


adder_full fa24_2(s23[3],c23[3],pr_and26[2],c24[3],s24[2]);


adder_full fa24_3(s23[4],c23[4],pr_and26[3],c24[4],s24[3]);


adder_full fa24_4(s23[5],c23[5],pr_and26[4],c24[5],s24[4]);


adder_full fa24_5(s23[6],c23[6],pr_and26[5],c24[6],s24[5]);


adder_full fa24_6(s23[7],c23[7],pr_and26[6],c24[7],s24[6]);


adder_full fa24_7(s23[8],c23[8],pr_and26[7],c24[8],s24[7]);


adder_full fa24_8(s23[9],c23[9],pr_and26[8],c24[9],s24[8]);


adder_full fa24_9(s23[10],c23[10],pr_and26[9],c24[10],s24[9]);


adder_full fa24_10(s23[11],c23[11],pr_and26[10],c24[11],s24[10]);


adder_full fa24_11(s23[12],c23[12],pr_and26[11],c24[12],s24[11]);


adder_full fa24_12(s23[13],c23[13],pr_and26[12],c24[13],s24[12]);


adder_full fa24_13(s23[14],c23[14],pr_and26[13],c24[14],s24[13]);


adder_full fa24_14(s23[15],c23[15],pr_and26[14],c24[15],s24[14]);


adder_full fa24_15(s23[16],c23[16],pr_and26[15],c24[16],s24[15]);


adder_full fa24_16(s23[17],c23[17],pr_and26[16],c24[17],s24[16]);


adder_full fa24_17(s23[18],c23[18],pr_and26[17],c24[18],s24[17]);


adder_full fa24_18(s23[19],c23[19],pr_and26[18],c24[19],s24[18]);


adder_full fa24_19(s23[20],c23[20],pr_and26[19],c24[20],s24[19]);


adder_full fa24_20(s23[21],c23[21],pr_and26[20],c24[21],s24[20]);


adder_full fa24_21(s23[22],c23[22],pr_and26[21],c24[22],s24[21]);


adder_full fa24_22(s23[23],c23[23],pr_and26[22],c24[23],s24[22]);


adder_full fa24_23(s23[24],c23[24],pr_and26[23],c24[24],s24[23]);


adder_full fa24_24(s23[25],c23[25],pr_and26[24],c24[25],s24[24]);


adder_full fa24_25(s23[26],c23[26],pr_and26[25],c24[26],s24[25]);


adder_full fa24_26(s23[27],c23[27],pr_and26[26],c24[27],s24[26]);


adder_full fa24_27(s23[28],c23[28],pr_and26[27],c24[28],s24[27]);


adder_full fa24_28(s23[29],c23[29],pr_and26[28],c24[29],s24[28]);


adder_full fa24_29(s23[30],c23[30],pr_and26[29],c24[30],s24[29]);


adder_full fa24_30(si[24],c23[31],pr_and26[30],c24[31],s24[30]);



//layer 25
adder_half ha25(s24[0],c24[0],c25[0],p[25]);


adder_full fa25_0(s24[1],c24[1],pr_and27[0],c25[1],s25[0]);


adder_full fa25_1(s24[2],c24[2],pr_and27[1],c25[2],s25[1]);


adder_full fa25_2(s24[3],c24[3],pr_and27[2],c25[3],s25[2]);


adder_full fa25_3(s24[4],c24[4],pr_and27[3],c25[4],s25[3]);


adder_full fa25_4(s24[5],c24[5],pr_and27[4],c25[5],s25[4]);


adder_full fa25_5(s24[6],c24[6],pr_and27[5],c25[6],s25[5]);


adder_full fa25_6(s24[7],c24[7],pr_and27[6],c25[7],s25[6]);


adder_full fa25_7(s24[8],c24[8],pr_and27[7],c25[8],s25[7]);


adder_full fa25_8(s24[9],c24[9],pr_and27[8],c25[9],s25[8]);


adder_full fa25_9(s24[10],c24[10],pr_and27[9],c25[10],s25[9]);


adder_full fa25_10(s24[11],c24[11],pr_and27[10],c25[11],s25[10]);


adder_full fa25_11(s24[12],c24[12],pr_and27[11],c25[12],s25[11]);


adder_full fa25_12(s24[13],c24[13],pr_and27[12],c25[13],s25[12]);


adder_full fa25_13(s24[14],c24[14],pr_and27[13],c25[14],s25[13]);


adder_full fa25_14(s24[15],c24[15],pr_and27[14],c25[15],s25[14]);


adder_full fa25_15(s24[16],c24[16],pr_and27[15],c25[16],s25[15]);


adder_full fa25_16(s24[17],c24[17],pr_and27[16],c25[17],s25[16]);


adder_full fa25_17(s24[18],c24[18],pr_and27[17],c25[18],s25[17]);


adder_full fa25_18(s24[19],c24[19],pr_and27[18],c25[19],s25[18]);


adder_full fa25_19(s24[20],c24[20],pr_and27[19],c25[20],s25[19]);


adder_full fa25_20(s24[21],c24[21],pr_and27[20],c25[21],s25[20]);


adder_full fa25_21(s24[22],c24[22],pr_and27[21],c25[22],s25[21]);


adder_full fa25_22(s24[23],c24[23],pr_and27[22],c25[23],s25[22]);


adder_full fa25_23(s24[24],c24[24],pr_and27[23],c25[24],s25[23]);


adder_full fa25_24(s24[25],c24[25],pr_and27[24],c25[25],s25[24]);


adder_full fa25_25(s24[26],c24[26],pr_and27[25],c25[26],s25[25]);


adder_full fa25_26(s24[27],c24[27],pr_and27[26],c25[27],s25[26]);


adder_full fa25_27(s24[28],c24[28],pr_and27[27],c25[28],s25[27]);


adder_full fa25_28(s24[29],c24[29],pr_and27[28],c25[29],s25[28]);


adder_full fa25_29(s24[30],c24[30],pr_and27[29],c25[30],s25[29]);


adder_full fa25_30(si[25],c24[31],pr_and27[30],c25[31],s25[30]);



//layer 26
adder_half ha26(s25[0],c25[0],c26[0],p[26]);


adder_full fa26_0(s25[1],c25[1],pr_and28[0],c26[1],s26[0]);


adder_full fa26_1(s25[2],c25[2],pr_and28[1],c26[2],s26[1]);


adder_full fa26_2(s25[3],c25[3],pr_and28[2],c26[3],s26[2]);


adder_full fa26_3(s25[4],c25[4],pr_and28[3],c26[4],s26[3]);


adder_full fa26_4(s25[5],c25[5],pr_and28[4],c26[5],s26[4]);


adder_full fa26_5(s25[6],c25[6],pr_and28[5],c26[6],s26[5]);


adder_full fa26_6(s25[7],c25[7],pr_and28[6],c26[7],s26[6]);


adder_full fa26_7(s25[8],c25[8],pr_and28[7],c26[8],s26[7]);


adder_full fa26_8(s25[9],c25[9],pr_and28[8],c26[9],s26[8]);


adder_full fa26_9(s25[10],c25[10],pr_and28[9],c26[10],s26[9]);


adder_full fa26_10(s25[11],c25[11],pr_and28[10],c26[11],s26[10]);


adder_full fa26_11(s25[12],c25[12],pr_and28[11],c26[12],s26[11]);


adder_full fa26_12(s25[13],c25[13],pr_and28[12],c26[13],s26[12]);


adder_full fa26_13(s25[14],c25[14],pr_and28[13],c26[14],s26[13]);


adder_full fa26_14(s25[15],c25[15],pr_and28[14],c26[15],s26[14]);


adder_full fa26_15(s25[16],c25[16],pr_and28[15],c26[16],s26[15]);


adder_full fa26_16(s25[17],c25[17],pr_and28[16],c26[17],s26[16]);


adder_full fa26_17(s25[18],c25[18],pr_and28[17],c26[18],s26[17]);


adder_full fa26_18(s25[19],c25[19],pr_and28[18],c26[19],s26[18]);


adder_full fa26_19(s25[20],c25[20],pr_and28[19],c26[20],s26[19]);


adder_full fa26_20(s25[21],c25[21],pr_and28[20],c26[21],s26[20]);


adder_full fa26_21(s25[22],c25[22],pr_and28[21],c26[22],s26[21]);


adder_full fa26_22(s25[23],c25[23],pr_and28[22],c26[23],s26[22]);


adder_full fa26_23(s25[24],c25[24],pr_and28[23],c26[24],s26[23]);


adder_full fa26_24(s25[25],c25[25],pr_and28[24],c26[25],s26[24]);


adder_full fa26_25(s25[26],c25[26],pr_and28[25],c26[26],s26[25]);


adder_full fa26_26(s25[27],c25[27],pr_and28[26],c26[27],s26[26]);


adder_full fa26_27(s25[28],c25[28],pr_and28[27],c26[28],s26[27]);


adder_full fa26_28(s25[29],c25[29],pr_and28[28],c26[29],s26[28]);


adder_full fa26_29(s25[30],c25[30],pr_and28[29],c26[30],s26[29]);


adder_full fa26_30(si[26],c25[31],pr_and28[30],c26[31],s26[30]);



//layer 27
adder_half ha27(s26[0],c26[0],c27[0],p[27]);


adder_full fa27_0(s26[1],c26[1],pr_and29[0],c27[1],s27[0]);


adder_full fa27_1(s26[2],c26[2],pr_and29[1],c27[2],s27[1]);


adder_full fa27_2(s26[3],c26[3],pr_and29[2],c27[3],s27[2]);


adder_full fa27_3(s26[4],c26[4],pr_and29[3],c27[4],s27[3]);


adder_full fa27_4(s26[5],c26[5],pr_and29[4],c27[5],s27[4]);


adder_full fa27_5(s26[6],c26[6],pr_and29[5],c27[6],s27[5]);


adder_full fa27_6(s26[7],c26[7],pr_and29[6],c27[7],s27[6]);


adder_full fa27_7(s26[8],c26[8],pr_and29[7],c27[8],s27[7]);


adder_full fa27_8(s26[9],c26[9],pr_and29[8],c27[9],s27[8]);


adder_full fa27_9(s26[10],c26[10],pr_and29[9],c27[10],s27[9]);


adder_full fa27_10(s26[11],c26[11],pr_and29[10],c27[11],s27[10]);


adder_full fa27_11(s26[12],c26[12],pr_and29[11],c27[12],s27[11]);


adder_full fa27_12(s26[13],c26[13],pr_and29[12],c27[13],s27[12]);


adder_full fa27_13(s26[14],c26[14],pr_and29[13],c27[14],s27[13]);


adder_full fa27_14(s26[15],c26[15],pr_and29[14],c27[15],s27[14]);


adder_full fa27_15(s26[16],c26[16],pr_and29[15],c27[16],s27[15]);


adder_full fa27_16(s26[17],c26[17],pr_and29[16],c27[17],s27[16]);


adder_full fa27_17(s26[18],c26[18],pr_and29[17],c27[18],s27[17]);


adder_full fa27_18(s26[19],c26[19],pr_and29[18],c27[19],s27[18]);


adder_full fa27_19(s26[20],c26[20],pr_and29[19],c27[20],s27[19]);


adder_full fa27_20(s26[21],c26[21],pr_and29[20],c27[21],s27[20]);


adder_full fa27_21(s26[22],c26[22],pr_and29[21],c27[22],s27[21]);


adder_full fa27_22(s26[23],c26[23],pr_and29[22],c27[23],s27[22]);


adder_full fa27_23(s26[24],c26[24],pr_and29[23],c27[24],s27[23]);


adder_full fa27_24(s26[25],c26[25],pr_and29[24],c27[25],s27[24]);


adder_full fa27_25(s26[26],c26[26],pr_and29[25],c27[26],s27[25]);


adder_full fa27_26(s26[27],c26[27],pr_and29[26],c27[27],s27[26]);


adder_full fa27_27(s26[28],c26[28],pr_and29[27],c27[28],s27[27]);


adder_full fa27_28(s26[29],c26[29],pr_and29[28],c27[29],s27[28]);


adder_full fa27_29(s26[30],c26[30],pr_and29[29],c27[30],s27[29]);


adder_full fa27_30(si[27],c26[31],pr_and29[30],c27[31],s27[30]);



//layer 28
adder_half ha28(s27[0],c27[0],c28[0],p[28]);


adder_full fa28_0(s27[1],c27[1],pr_and30[0],c28[1],s28[0]);


adder_full fa28_1(s27[2],c27[2],pr_and30[1],c28[2],s28[1]);


adder_full fa28_2(s27[3],c27[3],pr_and30[2],c28[3],s28[2]);


adder_full fa28_3(s27[4],c27[4],pr_and30[3],c28[4],s28[3]);


adder_full fa28_4(s27[5],c27[5],pr_and30[4],c28[5],s28[4]);


adder_full fa28_5(s27[6],c27[6],pr_and30[5],c28[6],s28[5]);


adder_full fa28_6(s27[7],c27[7],pr_and30[6],c28[7],s28[6]);


adder_full fa28_7(s27[8],c27[8],pr_and30[7],c28[8],s28[7]);


adder_full fa28_8(s27[9],c27[9],pr_and30[8],c28[9],s28[8]);


adder_full fa28_9(s27[10],c27[10],pr_and30[9],c28[10],s28[9]);


adder_full fa28_10(s27[11],c27[11],pr_and30[10],c28[11],s28[10]);


adder_full fa28_11(s27[12],c27[12],pr_and30[11],c28[12],s28[11]);


adder_full fa28_12(s27[13],c27[13],pr_and30[12],c28[13],s28[12]);


adder_full fa28_13(s27[14],c27[14],pr_and30[13],c28[14],s28[13]);


adder_full fa28_14(s27[15],c27[15],pr_and30[14],c28[15],s28[14]);


adder_full fa28_15(s27[16],c27[16],pr_and30[15],c28[16],s28[15]);


adder_full fa28_16(s27[17],c27[17],pr_and30[16],c28[17],s28[16]);


adder_full fa28_17(s27[18],c27[18],pr_and30[17],c28[18],s28[17]);


adder_full fa28_18(s27[19],c27[19],pr_and30[18],c28[19],s28[18]);


adder_full fa28_19(s27[20],c27[20],pr_and30[19],c28[20],s28[19]);


adder_full fa28_20(s27[21],c27[21],pr_and30[20],c28[21],s28[20]);


adder_full fa28_21(s27[22],c27[22],pr_and30[21],c28[22],s28[21]);


adder_full fa28_22(s27[23],c27[23],pr_and30[22],c28[23],s28[22]);


adder_full fa28_23(s27[24],c27[24],pr_and30[23],c28[24],s28[23]);


adder_full fa28_24(s27[25],c27[25],pr_and30[24],c28[25],s28[24]);


adder_full fa28_25(s27[26],c27[26],pr_and30[25],c28[26],s28[25]);


adder_full fa28_26(s27[27],c27[27],pr_and30[26],c28[27],s28[26]);


adder_full fa28_27(s27[28],c27[28],pr_and30[27],c28[28],s28[27]);


adder_full fa28_28(s27[29],c27[29],pr_and30[28],c28[29],s28[28]);


adder_full fa28_29(s27[30],c27[30],pr_and30[29],c28[30],s28[29]);


adder_full fa28_30(si[28],c27[31],pr_and30[30],c28[31],s28[30]);



//layer 29
adder_half ha29(s28[0],c28[0],c29[0],p[29]);


adder_full fa29_0(s28[1],c28[1],pr_and31[0],c29[1],s29[0]);


adder_full fa29_1(s28[2],c28[2],pr_and31[1],c29[2],s29[1]);


adder_full fa29_2(s28[3],c28[3],pr_and31[2],c29[3],s29[2]);


adder_full fa29_3(s28[4],c28[4],pr_and31[3],c29[4],s29[3]);


adder_full fa29_4(s28[5],c28[5],pr_and31[4],c29[5],s29[4]);


adder_full fa29_5(s28[6],c28[6],pr_and31[5],c29[6],s29[5]);


adder_full fa29_6(s28[7],c28[7],pr_and31[6],c29[7],s29[6]);


adder_full fa29_7(s28[8],c28[8],pr_and31[7],c29[8],s29[7]);


adder_full fa29_8(s28[9],c28[9],pr_and31[8],c29[9],s29[8]);


adder_full fa29_9(s28[10],c28[10],pr_and31[9],c29[10],s29[9]);


adder_full fa29_10(s28[11],c28[11],pr_and31[10],c29[11],s29[10]);


adder_full fa29_11(s28[12],c28[12],pr_and31[11],c29[12],s29[11]);


adder_full fa29_12(s28[13],c28[13],pr_and31[12],c29[13],s29[12]);


adder_full fa29_13(s28[14],c28[14],pr_and31[13],c29[14],s29[13]);


adder_full fa29_14(s28[15],c28[15],pr_and31[14],c29[15],s29[14]);


adder_full fa29_15(s28[16],c28[16],pr_and31[15],c29[16],s29[15]);


adder_full fa29_16(s28[17],c28[17],pr_and31[16],c29[17],s29[16]);


adder_full fa29_17(s28[18],c28[18],pr_and31[17],c29[18],s29[17]);


adder_full fa29_18(s28[19],c28[19],pr_and31[18],c29[19],s29[18]);


adder_full fa29_19(s28[20],c28[20],pr_and31[19],c29[20],s29[19]);


adder_full fa29_20(s28[21],c28[21],pr_and31[20],c29[21],s29[20]);


adder_full fa29_21(s28[22],c28[22],pr_and31[21],c29[22],s29[21]);


adder_full fa29_22(s28[23],c28[23],pr_and31[22],c29[23],s29[22]);


adder_full fa29_23(s28[24],c28[24],pr_and31[23],c29[24],s29[23]);


adder_full fa29_24(s28[25],c28[25],pr_and31[24],c29[25],s29[24]);


adder_full fa29_25(s28[26],c28[26],pr_and31[25],c29[26],s29[25]);


adder_full fa29_26(s28[27],c28[27],pr_and31[26],c29[27],s29[26]);


adder_full fa29_27(s28[28],c28[28],pr_and31[27],c29[28],s29[27]);


adder_full fa29_28(s28[29],c28[29],pr_and31[28],c29[29],s29[28]);


adder_full fa29_29(s28[30],c28[30],pr_and31[29],c29[30],s29[29]);


adder_full fa29_30(si[29],c28[31],pr_and31[30],c29[31],s29[30]);



//layer 30
adder_half ha30(s29[0],c29[0],c30[0],p[30]);


adder_full fa30_0(s29[1],c29[1],pr_and32[0],c30[1],s30[0]);


adder_full fa30_1(s29[2],c29[2],pr_and32[1],c30[2],s30[1]);


adder_full fa30_2(s29[3],c29[3],pr_and32[2],c30[3],s30[2]);


adder_full fa30_3(s29[4],c29[4],pr_and32[3],c30[4],s30[3]);


adder_full fa30_4(s29[5],c29[5],pr_and32[4],c30[5],s30[4]);


adder_full fa30_5(s29[6],c29[6],pr_and32[5],c30[6],s30[5]);


adder_full fa30_6(s29[7],c29[7],pr_and32[6],c30[7],s30[6]);


adder_full fa30_7(s29[8],c29[8],pr_and32[7],c30[8],s30[7]);


adder_full fa30_8(s29[9],c29[9],pr_and32[8],c30[9],s30[8]);


adder_full fa30_9(s29[10],c29[10],pr_and32[9],c30[10],s30[9]);


adder_full fa30_10(s29[11],c29[11],pr_and32[10],c30[11],s30[10]);


adder_full fa30_11(s29[12],c29[12],pr_and32[11],c30[12],s30[11]);


adder_full fa30_12(s29[13],c29[13],pr_and32[12],c30[13],s30[12]);


adder_full fa30_13(s29[14],c29[14],pr_and32[13],c30[14],s30[13]);


adder_full fa30_14(s29[15],c29[15],pr_and32[14],c30[15],s30[14]);


adder_full fa30_15(s29[16],c29[16],pr_and32[15],c30[16],s30[15]);


adder_full fa30_16(s29[17],c29[17],pr_and32[16],c30[17],s30[16]);


adder_full fa30_17(s29[18],c29[18],pr_and32[17],c30[18],s30[17]);


adder_full fa30_18(s29[19],c29[19],pr_and32[18],c30[19],s30[18]);


adder_full fa30_19(s29[20],c29[20],pr_and32[19],c30[20],s30[19]);


adder_full fa30_20(s29[21],c29[21],pr_and32[20],c30[21],s30[20]);


adder_full fa30_21(s29[22],c29[22],pr_and32[21],c30[22],s30[21]);


adder_full fa30_22(s29[23],c29[23],pr_and32[22],c30[23],s30[22]);


adder_full fa30_23(s29[24],c29[24],pr_and32[23],c30[24],s30[23]);


adder_full fa30_24(s29[25],c29[25],pr_and32[24],c30[25],s30[24]);


adder_full fa30_25(s29[26],c29[26],pr_and32[25],c30[26],s30[25]);


adder_full fa30_26(s29[27],c29[27],pr_and32[26],c30[27],s30[26]);


adder_full fa30_27(s29[28],c29[28],pr_and32[27],c30[28],s30[27]);


adder_full fa30_28(s29[29],c29[29],pr_and32[28],c30[29],s30[28]);


adder_full fa30_29(s29[30],c29[30],pr_and32[29],c30[30],s30[29]);


adder_full fa30_30(si[30],c29[31],pr_and32[30],c30[31],s30[30]);



//last layer
adder_full fad31_30(s30[0],c30[0],b[31],c31[0],p[31]);


adder_full fad31_31(s30[1],c30[1],c31[0],c31[1],p[32]);


adder_full fad31_32(s30[2],c30[2],c31[1],c31[2],p[33]);


adder_full fad31_33(s30[3],c30[3],c31[2],c31[3],p[34]);


adder_full fad31_34(s30[4],c30[4],c31[3],c31[4],p[35]);


adder_full fad31_35(s30[5],c30[5],c31[4],c31[5],p[36]);


adder_full fad31_36(s30[6],c30[6],c31[5],c31[6],p[37]);


adder_full fad31_37(s30[7],c30[7],c31[6],c31[7],p[38]);


adder_full fad31_38(s30[8],c30[8],c31[7],c31[8],p[39]);


adder_full fad31_39(s30[9],c30[9],c31[8],c31[9],p[40]);


adder_full fad31_40(s30[10],c30[10],c31[9],c31[10],p[41]);


adder_full fad31_41(s30[11],c30[11],c31[10],c31[11],p[42]);


adder_full fad31_42(s30[12],c30[12],c31[11],c31[12],p[43]);


adder_full fad31_43(s30[13],c30[13],c31[12],c31[13],p[44]);


adder_full fad31_44(s30[14],c30[14],c31[13],c31[14],p[45]);


adder_full fad31_45(s30[15],c30[15],c31[14],c31[15],p[46]);


adder_full fad31_46(s30[16],c30[16],c31[15],c31[16],p[47]);


adder_full fad31_47(s30[17],c30[17],c31[16],c31[17],p[48]);


adder_full fad31_48(s30[18],c30[18],c31[17],c31[18],p[49]);


adder_full fad31_49(s30[19],c30[19],c31[18],c31[19],p[50]);


adder_full fad31_50(s30[20],c30[20],c31[19],c31[20],p[51]);


adder_full fad31_51(s30[21],c30[21],c31[20],c31[21],p[52]);


adder_full fad31_52(s30[22],c30[22],c31[21],c31[22],p[53]);


adder_full fad31_53(s30[23],c30[23],c31[22],c31[23],p[54]);


adder_full fad31_54(s30[24],c30[24],c31[23],c31[24],p[55]);


adder_full fad31_55(s30[25],c30[25],c31[24],c31[25],p[56]);


adder_full fad31_56(s30[26],c30[26],c31[25],c31[26],p[57]);


adder_full fad31_57(s30[27],c30[27],c31[26],c31[27],p[58]);


adder_full fad31_58(s30[28],c30[28],c31[27],c31[28],p[59]);


adder_full fad31_59(s30[29],c30[29],c31[28],c31[29],p[60]);


adder_full fad31_60(s30[30],c30[30],c31[29],c31[30],p[61]);


adder_full fad31_61(si[31],c30[31],c31[30],c31[31],p[62]);
adder_half ha32(c31[31],1'b1,c,p[63]);
assign p[0]=pr_and1[0];

endmodule